--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity Losing_Sound is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(14 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end Losing_Sound;

architecture arch of Losing_Sound is
constant array_size 			: integer := 26574 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal sin_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
  sintable_proc: process(resetN, CLK)
    constant sin_table : table_type := (
---start 0 v

X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"007D",
X"FF06",
X"FE0C",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"0177",
X"01F4",
X"0271",
X"0271",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"007D",
X"FF06",
X"FE0C",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"007D",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0177",
X"0000",
X"FE89",
X"FD12",
X"FC18",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FD8F",
X"FE89",
X"0000",
X"007D",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"00FA",
X"007D",
X"007D",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"02EE",
X"0271",
X"00FA",
X"FF83",
X"FD8F",
X"FC95",
X"FB9B",
X"FB1E",
X"FB1E",
X"FC18",
X"FD12",
X"FE0C",
X"FF83",
X"007D",
X"0177",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"00FA",
X"007D",
X"0000",
X"0000",
X"00FA",
X"0177",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"007D",
X"FE89",
X"FC95",
X"FB9B",
X"FAA1",
X"FAA1",
X"FB9B",
X"FC95",
X"FD8F",
X"FF06",
X"007D",
X"0177",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0177",
X"007D",
X"0000",
X"0000",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"02EE",
X"0177",
X"FF06",
X"FD12",
X"FB9B",
X"FAA1",
X"FAA1",
X"FAA1",
X"FB9B",
X"FD12",
X"FE89",
X"0000",
X"0177",
X"0271",
X"02EE",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"00FA",
X"0000",
X"0000",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"036B",
X"01F4",
X"0000",
X"FE0C",
X"FC18",
X"FB1E",
X"FAA1",
X"FAA1",
X"FB1E",
X"FC95",
X"FD8F",
X"FF06",
X"007D",
X"01F4",
X"02EE",
X"036B",
X"036B",
X"02EE",
X"0271",
X"0177",
X"007D",
X"0000",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"02EE",
X"02EE",
X"0271",
X"0177",
X"0000",
X"FE0C",
X"FC18",
X"FB1E",
X"FA24",
X"FAA1",
X"FB9B",
X"FC95",
X"FE0C",
X"FF83",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"036B",
X"02EE",
X"01F4",
X"00FA",
X"007D",
X"0000",
X"0000",
X"007D",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0177",
X"00FA",
X"FF83",
X"FE89",
X"FD12",
X"FC18",
X"FB9B",
X"FB9B",
X"FC18",
X"FD12",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"0271",
X"01F4",
X"00FA",
X"0000",
X"FE89",
X"FD8F",
X"FC95",
X"FB9B",
X"FB9B",
X"FC18",
X"FD12",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"02EE",
X"0271",
X"0177",
X"0000",
X"FE89",
X"FD12",
X"FC18",
X"FB9B",
X"FB9B",
X"FC95",
X"FD8F",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"01F4",
X"0000",
X"FE89",
X"FD12",
X"FC18",
X"FB1E",
X"FB1E",
X"FB9B",
X"FD12",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"00FA",
X"0177",
X"02EE",
X"036B",
X"036B",
X"0271",
X"00FA",
X"FF83",
X"FD8F",
X"FC18",
X"FB1E",
X"FAA1",
X"FAA1",
X"FC18",
X"FD8F",
X"FF06",
X"0000",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"0177",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"007D",
X"01F4",
X"02EE",
X"03E8",
X"03E8",
X"0271",
X"00FA",
X"FF06",
X"FD8F",
X"FC18",
X"FAA1",
X"FA24",
X"FAA1",
X"FB9B",
X"FD12",
X"FE89",
X"0000",
X"0177",
X"0271",
X"02EE",
X"036B",
X"02EE",
X"0271",
X"0177",
X"007D",
X"FF83",
X"FF06",
X"FF06",
X"0000",
X"0177",
X"02EE",
X"03E8",
X"03E8",
X"036B",
X"01F4",
X"0000",
X"FE89",
X"FD12",
X"FB9B",
X"FAA1",
X"FAA1",
X"FB1E",
X"FC95",
X"FE0C",
X"FF83",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"00FA",
X"FF83",
X"FF06",
X"FE89",
X"FF06",
X"007D",
X"01F4",
X"036B",
X"03E8",
X"036B",
X"0271",
X"00FA",
X"FF06",
X"FD8F",
X"FC18",
X"FB1E",
X"FAA1",
X"FB1E",
X"FC95",
X"FE0C",
X"FF06",
X"007D",
X"0177",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"FF83",
X"007D",
X"01F4",
X"02EE",
X"036B",
X"02EE",
X"01F4",
X"007D",
X"FE89",
X"FC95",
X"FB9B",
X"FAA1",
X"FAA1",
X"FB9B",
X"FD12",
X"FE89",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"00FA",
X"0000",
X"FF83",
X"0000",
X"007D",
X"01F4",
X"02EE",
X"036B",
X"02EE",
X"01F4",
X"007D",
X"FE89",
X"FC95",
X"FB1E",
X"FAA1",
X"FAA1",
X"FB1E",
X"FC95",
X"FE0C",
X"FF83",
X"007D",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"0271",
X"0271",
X"0177",
X"007D",
X"0000",
X"0000",
X"007D",
X"01F4",
X"036B",
X"03E8",
X"03E8",
X"0271",
X"007D",
X"FE89",
X"FC95",
X"FAA1",
X"F9A7",
X"F92A",
X"FA24",
X"FB9B",
X"FD8F",
X"FF06",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"03E8",
X"036B",
X"02EE",
X"01F4",
X"007D",
X"0000",
X"FF83",
X"0000",
X"00FA",
X"0271",
X"03E8",
X"03E8",
X"02EE",
X"0177",
X"FF83",
X"FD8F",
X"FB9B",
X"FA24",
X"F92A",
X"F92A",
X"FAA1",
X"FC18",
X"FE0C",
X"FF83",
X"0177",
X"02EE",
X"03E8",
X"0465",
X"0465",
X"036B",
X"02EE",
X"0177",
X"0000",
X"FF06",
X"FF06",
X"FF83",
X"00FA",
X"0271",
X"03E8",
X"036B",
X"0271",
X"00FA",
X"FF83",
X"FD8F",
X"FC18",
X"FAA1",
X"F9A7",
X"F9A7",
X"FAA1",
X"FC95",
X"FE0C",
X"0000",
X"0177",
X"0271",
X"03E8",
X"0465",
X"03E8",
X"036B",
X"0271",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"FF83",
X"00FA",
X"0271",
X"036B",
X"036B",
X"0271",
X"00FA",
X"FF83",
X"FE0C",
X"FC18",
X"FB1E",
X"FA24",
X"FAA1",
X"FB9B",
X"FD12",
X"FE89",
X"0000",
X"0177",
X"0271",
X"036B",
X"036B",
X"036B",
X"02EE",
X"01F4",
X"00FA",
X"0000",
X"FF83",
X"FF83",
X"007D",
X"0177",
X"02EE",
X"036B",
X"02EE",
X"01F4",
X"007D",
X"FE89",
X"FD12",
X"FB9B",
X"FA24",
X"FA24",
X"FB1E",
X"FC18",
X"FE0C",
X"FF83",
X"007D",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0177",
X"007D",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"036B",
X"03E8",
X"036B",
X"01F4",
X"0000",
X"FE0C",
X"FC18",
X"FA24",
X"F9A7",
X"F9A7",
X"FAA1",
X"FC18",
X"FE0C",
X"FF83",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"036B",
X"02EE",
X"0271",
X"0177",
X"00FA",
X"007D",
X"007D",
X"00FA",
X"0271",
X"03E8",
X"04E2",
X"03E8",
X"0271",
X"0000",
X"FD8F",
X"FB1E",
X"F92A",
X"F830",
X"F830",
X"F9A7",
X"FB1E",
X"FD8F",
X"FF06",
X"00FA",
X"0271",
X"036B",
X"03E8",
X"0465",
X"03E8",
X"02EE",
X"01F4",
X"00FA",
X"0000",
X"007D",
X"0177",
X"0271",
X"03E8",
X"04E2",
X"0465",
X"02EE",
X"007D",
X"FE0C",
X"FB9B",
X"F9A7",
X"F830",
X"F7B3",
X"F8AD",
X"FAA1",
X"FC95",
X"FE89",
X"0000",
X"01F4",
X"036B",
X"0465",
X"04E2",
X"0465",
X"03E8",
X"0271",
X"00FA",
X"0000",
X"0000",
X"00FA",
X"01F4",
X"036B",
X"0465",
X"0465",
X"02EE",
X"00FA",
X"FE89",
X"FC95",
X"FAA1",
X"F92A",
X"F830",
X"F830",
X"F9A7",
X"FB9B",
X"FD8F",
X"FF06",
X"00FA",
X"0271",
X"03E8",
X"04E2",
X"04E2",
X"03E8",
X"02EE",
X"0177",
X"007D",
X"0000",
X"007D",
X"0177",
X"0271",
X"03E8",
X"0465",
X"03E8",
X"01F4",
X"0000",
X"FD8F",
X"FB9B",
X"FA24",
X"F92A",
X"F830",
X"F92A",
X"FAA1",
X"FC95",
X"FE89",
X"007D",
X"01F4",
X"036B",
X"0465",
X"04E2",
X"03E8",
X"02EE",
X"01F4",
X"007D",
X"0000",
X"0000",
X"00FA",
X"01F4",
X"03E8",
X"0465",
X"0465",
X"02EE",
X"007D",
X"FE0C",
X"FC18",
X"FA24",
X"F8AD",
X"F7B3",
X"F830",
X"FA24",
X"FC95",
X"FE89",
X"007D",
X"01F4",
X"036B",
X"0465",
X"04E2",
X"03E8",
X"036B",
X"01F4",
X"00FA",
X"007D",
X"007D",
X"0177",
X"0271",
X"03E8",
X"04E2",
X"0465",
X"02EE",
X"007D",
X"FE0C",
X"FB9B",
X"F92A",
X"F7B3",
X"F6B9",
X"F7B3",
X"F9A7",
X"FC18",
X"FE89",
X"007D",
X"02EE",
X"0465",
X"055F",
X"055F",
X"04E2",
X"03E8",
X"0271",
X"00FA",
X"007D",
X"007D",
X"0177",
X"02EE",
X"0465",
X"055F",
X"04E2",
X"02EE",
X"0000",
X"FD12",
X"FA24",
X"F830",
X"F63C",
X"F542",
X"F6B9",
X"F92A",
X"FC18",
X"FE89",
X"0177",
X"036B",
X"04E2",
X"05DC",
X"05DC",
X"055F",
X"0465",
X"02EE",
X"0177",
X"007D",
X"00FA",
X"01F4",
X"036B",
X"04E2",
X"055F",
X"04E2",
X"02EE",
X"0000",
X"FC95",
X"F9A7",
X"F736",
X"F542",
X"F448",
X"F5BF",
X"F8AD",
X"FB9B",
X"FE0C",
X"00FA",
X"03E8",
X"05DC",
X"06D6",
X"06D6",
X"05DC",
X"04E2",
X"036B",
X"01F4",
X"00FA",
X"00FA",
X"0271",
X"03E8",
X"04E2",
X"055F",
X"0465",
X"0271",
X"0000",
X"FC95",
X"F92A",
X"F736",
X"F542",
X"F448",
X"F542",
X"F7B3",
X"FB1E",
X"FE0C",
X"00FA",
X"036B",
X"05DC",
X"06D6",
X"0753",
X"06D6",
X"055F",
X"03E8",
X"0271",
X"00FA",
X"00FA",
X"01F4",
X"036B",
X"04E2",
X"055F",
X"0465",
X"0271",
X"0000",
X"FC95",
X"F9A7",
X"F736",
X"F5BF",
X"F4C5",
X"F542",
X"F7B3",
X"FAA1",
X"FD8F",
X"0000",
X"02EE",
X"055F",
X"06D6",
X"0753",
X"06D6",
X"05DC",
X"0465",
X"02EE",
X"0177",
X"00FA",
X"01F4",
X"02EE",
X"03E8",
X"04E2",
X"04E2",
X"036B",
X"007D",
X"FD12",
X"F9A7",
X"F736",
X"F5BF",
X"F448",
X"F4C5",
X"F736",
X"FAA1",
X"FD8F",
X"007D",
X"036B",
X"055F",
X"06D6",
X"0753",
X"06D6",
X"05DC",
X"0465",
X"0271",
X"0177",
X"00FA",
X"01F4",
X"02EE",
X"0465",
X"055F",
X"055F",
X"036B",
X"007D",
X"FD12",
X"F9A7",
X"F6B9",
X"F448",
X"F2D1",
X"F448",
X"F736",
X"FAA1",
X"FE0C",
X"00FA",
X"03E8",
X"0659",
X"07D0",
X"07D0",
X"06D6",
X"05DC",
X"0465",
X"0271",
X"00FA",
X"00FA",
X"01F4",
X"036B",
X"055F",
X"0659",
X"05DC",
X"03E8",
X"007D",
X"FC18",
X"F8AD",
X"F542",
X"F2D1",
X"F1D7",
X"F34E",
X"F6B9",
X"FAA1",
X"FE0C",
X"01F4",
X"04E2",
X"0753",
X"08CA",
X"08CA",
X"07D0",
X"05DC",
X"03E8",
X"01F4",
X"007D",
X"007D",
X"0177",
X"036B",
X"055F",
X"06D6",
X"0659",
X"0465",
X"007D",
X"FC95",
X"F830",
X"F4C5",
X"F1D7",
X"F15A",
X"F2D1",
X"F63C",
X"FA24",
X"FE0C",
X"01F4",
X"055F",
X"084D",
X"0947",
X"0947",
X"07D0",
X"0659",
X"03E8",
X"01F4",
X"007D",
X"0000",
X"00FA",
X"02EE",
X"04E2",
X"0659",
X"0659",
X"0465",
X"0177",
X"FD12",
X"F8AD",
X"F542",
X"F1D7",
X"F0DD",
X"F254",
X"F542",
X"F92A",
X"FD8F",
X"0177",
X"055F",
X"07D0",
X"09C4",
X"09C4",
X"08CA",
X"06D6",
X"0465",
X"01F4",
X"007D",
X"0000",
X"007D",
X"0271",
X"04E2",
X"0659",
X"0659",
X"04E2",
X"0177",
X"FD12",
X"F8AD",
X"F542",
X"F254",
X"F15A",
X"F254",
X"F542",
X"F92A",
X"FD8F",
X"0177",
X"055F",
X"07D0",
X"09C4",
X"09C4",
X"08CA",
X"06D6",
X"0465",
X"01F4",
X"0000",
X"FF83",
X"007D",
X"01F4",
X"04E2",
X"06D6",
X"0753",
X"05DC",
X"0271",
X"FD8F",
X"F92A",
X"F4C5",
X"F1D7",
X"F060",
X"F1D7",
X"F4C5",
X"F92A",
X"FD8F",
X"0177",
X"055F",
X"084D",
X"09C4",
X"09C4",
X"08CA",
X"06D6",
X"0465",
X"0177",
X"0000",
X"FF83",
X"007D",
X"01F4",
X"04E2",
X"06D6",
X"07D0",
X"06D6",
X"036B",
X"FE0C",
X"F92A",
X"F448",
X"F0DD",
X"EF66",
X"F0DD",
X"F448",
X"F830",
X"FD12",
X"0177",
X"055F",
X"084D",
X"09C4",
X"09C4",
X"08CA",
X"0753",
X"0465",
X"01F4",
X"0000",
X"FF83",
X"007D",
X"0271",
X"04E2",
X"0753",
X"08CA",
X"0753",
X"03E8",
X"FE89",
X"F8AD",
X"F3CB",
X"EFE3",
X"EEE9",
X"F060",
X"F3CB",
X"F830",
X"FC95",
X"0177",
X"055F",
X"084D",
X"09C4",
X"0A41",
X"0947",
X"0753",
X"04E2",
X"01F4",
X"0000",
X"FF83",
X"007D",
X"02EE",
X"055F",
X"07D0",
X"0947",
X"07D0",
X"03E8",
X"FE89",
X"F830",
X"F2D1",
X"EEE9",
X"EDEF",
X"EF66",
X"F34E",
X"F7B3",
X"FC95",
X"0177",
X"05DC",
X"08CA",
X"0A41",
X"0ABE",
X"09C4",
X"07D0",
X"04E2",
X"01F4",
X"0000",
X"FF06",
X"0000",
X"0271",
X"055F",
X"084D",
X"09C4",
X"084D",
X"0465",
X"FE89",
X"F8AD",
X"F2D1",
X"EEE9",
X"ED72",
X"EF66",
X"F2D1",
X"F736",
X"FC18",
X"00FA",
X"055F",
X"08CA",
X"0A41",
X"0ABE",
X"09C4",
X"07D0",
X"055F",
X"0271",
X"0000",
X"FF83",
X"0000",
X"01F4",
X"04E2",
X"07D0",
X"0947",
X"084D",
X"04E2",
X"FF06",
X"F8AD",
X"F2D1",
X"EEE9",
X"ED72",
X"EF66",
X"F2D1",
X"F7B3",
X"FD12",
X"0177",
X"05DC",
X"0947",
X"0A41",
X"0A41",
X"0947",
X"07D0",
X"04E2",
X"01F4",
X"0000",
X"FF06",
X"FF83",
X"01F4",
X"04E2",
X"07D0",
X"09C4",
X"08CA",
X"055F",
X"FF83",
X"F92A",
X"F254",
X"EDEF",
X"EC78",
X"EE6C",
X"F2D1",
X"F7B3",
X"FD12",
X"01F4",
X"0659",
X"0947",
X"0A41",
X"0A41",
X"0947",
X"0753",
X"04E2",
X"01F4",
X"0000",
X"FF06",
X"FF83",
X"01F4",
X"04E2",
X"07D0",
X"0A41",
X"0A41",
X"06D6",
X"00FA",
X"F9A7",
X"F254",
X"ED72",
X"EB7E",
X"ED72",
X"F1D7",
X"F6B9",
X"FC95",
X"01F4",
X"0659",
X"0947",
X"0ABE",
X"0ABE",
X"09C4",
X"084D",
X"055F",
X"01F4",
X"FF83",
X"FE89",
X"FF06",
X"0177",
X"04E2",
X"084D",
X"0ABE",
X"0ABE",
X"07D0",
X"0177",
X"FA24",
X"F254",
X"EC78",
X"EA84",
X"EC78",
X"F0DD",
X"F63C",
X"FC18",
X"0177",
X"0659",
X"09C4",
X"0B3B",
X"0B3B",
X"0A41",
X"084D",
X"055F",
X"0177",
X"FF06",
X"FE89",
X"FF06",
X"00FA",
X"0465",
X"084D",
X"0B3B",
X"0C35",
X"0947",
X"036B",
X"FB1E",
X"F1D7",
X"EB7E",
X"E90D",
X"EB01",
X"EF66",
X"F4C5",
X"FB1E",
X"0177",
X"06D6",
X"0A41",
X"0BB8",
X"0BB8",
X"0ABE",
X"08CA",
X"055F",
X"01F4",
X"FF83",
X"FF06",
X"FF06",
X"00FA",
X"03E8",
X"07D0",
X"0ABE",
X"0BB8",
X"09C4",
X"036B",
X"FB1E",
X"F1D7",
X"EB7E",
X"E90D",
X"EA84",
X"EF66",
X"F542",
X"FB9B",
X"0177",
X"06D6",
X"0A41",
X"0BB8",
X"0BB8",
X"0ABE",
X"0947",
X"05DC",
X"0271",
X"0000",
X"FF06",
X"FF06",
X"007D",
X"03E8",
X"07D0",
X"0BB8",
X"0D2F",
X"0ABE",
X"03E8",
X"FB1E",
X"F1D7",
X"EB01",
X"E813",
X"EA07",
X"EE6C",
X"F3CB",
X"FAA1",
X"00FA",
X"0659",
X"0A41",
X"0BB8",
X"0BB8",
X"0B3B",
X"09C4",
X"0659",
X"0271",
X"FF83",
X"FE89",
X"FE89",
X"007D",
X"036B",
X"07D0",
X"0B3B",
X"0CB2",
X"0ABE",
X"055F",
X"FC95",
X"F34E",
X"EBFB",
X"E890",
X"EA07",
X"EE6C",
X"F3CB",
X"FA24",
X"0000",
X"05DC",
X"0947",
X"0B3B",
X"0BB8",
X"0B3B",
X"0947",
X"0659",
X"02EE",
X"0000",
X"FE89",
X"FE89",
X"0000",
X"02EE",
X"06D6",
X"0ABE",
X"0CB2",
X"0BB8",
X"0659",
X"FE0C",
X"F448",
X"EBFB",
X"E890",
X"EA07",
X"EE6C",
X"F3CB",
X"F9A7",
X"0000",
X"05DC",
X"0947",
X"0ABE",
X"0ABE",
X"0A41",
X"08CA",
X"0659",
X"02EE",
X"007D",
X"FF06",
X"FE89",
X"0000",
X"0271",
X"0659",
X"0ABE",
X"0DAC",
X"0CB2",
X"0753",
X"FE89",
X"F4C5",
X"EBFB",
X"E813",
X"E90D",
X"ED72",
X"F34E",
X"F9A7",
X"0000",
X"05DC",
X"0947",
X"0ABE",
X"0ABE",
X"0ABE",
X"0947",
X"0659",
X"02EE",
X"0000",
X"FE89",
X"FE0C",
X"FF06",
X"0271",
X"06D6",
X"0B3B",
X"0E29",
X"0DAC",
X"084D",
X"FF06",
X"F4C5",
X"EB7E",
X"E719",
X"E890",
X"ECF5",
X"F254",
X"F92A",
X"0000",
X"05DC",
X"0947",
X"0B3B",
X"0B3B",
X"0ABE",
X"09C4",
X"06D6",
X"036B",
X"007D",
X"FE89",
X"FE0C",
X"FF06",
X"01F4",
X"0659",
X"0BB8",
X"0F23",
X"0EA6",
X"0947",
X"FF06",
X"F448",
X"EA84",
X"E69C",
X"E813",
X"EC78",
X"F1D7",
X"F8AD",
X"FF83",
X"05DC",
X"09C4",
X"0B3B",
X"0BB8",
X"0B3B",
X"09C4",
X"06D6",
X"036B",
X"0000",
X"FE89",
X"FE0C",
X"FF83",
X"0271",
X"06D6",
X"0C35",
X"101D",
X"0F23",
X"0947",
X"FE89",
X"F2D1",
X"E98A",
X"E5A2",
X"E719",
X"EB7E",
X"F1D7",
X"F92A",
X"007D",
X"0659",
X"0A41",
X"0BB8",
X"0C35",
X"0BB8",
X"0A41",
X"0753",
X"036B",
X"007D",
X"FE89",
X"FE0C",
X"FF06",
X"01F4",
X"06D6",
X"0C35",
X"101D",
X"0F23",
X"08CA",
X"FE0C",
X"F2D1",
X"E90D",
X"E4A8",
X"E69C",
X"EB7E",
X"F15A",
X"F8AD",
X"007D",
X"06D6",
X"0ABE",
X"0C35",
X"0CB2",
X"0CB2",
X"0ABE",
X"0753",
X"036B",
X"0000",
X"FD8F",
X"FD8F",
X"FE89",
X"01F4",
X"0659",
X"0BB8",
X"0FA0",
X"0F23",
X"09C4",
X"FF83",
X"F3CB",
X"E98A",
X"E525",
X"E69C",
X"EA84",
X"F060",
X"F7B3",
X"FF83",
X"05DC",
X"0A41",
X"0CB2",
X"0D2F",
X"0D2F",
X"0B3B",
X"07D0",
X"03E8",
X"0000",
X"FE0C",
X"FD8F",
X"FF06",
X"01F4",
X"0659",
X"0BB8",
X"101D",
X"0FA0",
X"0A41",
X"0000",
X"F3CB",
X"E90D",
X"E42B",
X"E5A2",
X"E98A",
X"EFE3",
X"F736",
X"FF83",
X"06D6",
X"0B3B",
X"0DAC",
X"0DAC",
X"0D2F",
X"0B3B",
X"0753",
X"036B",
X"0000",
X"FD8F",
X"FD8F",
X"FF06",
X"01F4",
X"0659",
X"0C35",
X"101D",
X"0FA0",
X"0ABE",
X"00FA",
X"F448",
X"E90D",
X"E42B",
X"E5A2",
X"EA07",
X"EF66",
X"F6B9",
X"FF06",
X"05DC",
X"0ABE",
X"0D2F",
X"0DAC",
X"0D2F",
X"0B3B",
X"0753",
X"02EE",
X"0000",
X"FE0C",
X"FE0C",
X"FF83",
X"02EE",
X"06D6",
X"0BB8",
X"0FA0",
X"0FA0",
X"0B3B",
X"01F4",
X"F4C5",
X"E90D",
X"E4A8",
X"E61F",
X"E98A",
X"EEE9",
X"F63C",
X"FE89",
X"055F",
X"0ABE",
X"0D2F",
X"0DAC",
X"0D2F",
X"0ABE",
X"06D6",
X"02EE",
X"0000",
X"FE0C",
X"FE0C",
X"0000",
X"0271",
X"0659",
X"0B3B",
X"0FA0",
X"109A",
X"0C35",
X"0271",
X"F4C5",
X"E813",
X"E3AE",
X"E525",
X"E90D",
X"EE6C",
X"F63C",
X"FF06",
X"0659",
X"0B3B",
X"0DAC",
X"0DAC",
X"0CB2",
X"0ABE",
X"0753",
X"02EE",
X"FF83",
X"FE0C",
X"FE0C",
X"FF06",
X"01F4",
X"0659",
X"0C35",
X"1117",
X"1211",
X"0D2F",
X"0271",
X"F448",
X"E813",
X"E331",
X"E4A8",
X"E796",
X"ED72",
X"F5BF",
X"FE89",
X"06D6",
X"0C35",
X"0E29",
X"0EA6",
X"0DAC",
X"0ABE",
X"06D6",
X"0271",
X"FE89",
X"FC95",
X"FD12",
X"FE89",
X"01F4",
X"06D6",
X"0D2F",
X"1211",
X"130B",
X"0E29",
X"02EE",
X"F448",
X"E796",
X"E2B4",
X"E3AE",
X"E69C",
X"EC78",
X"F5BF",
X"FF83",
X"0753",
X"0D2F",
X"0FA0",
X"0FA0",
X"0E29",
X"0ABE",
X"0659",
X"0177",
X"FD8F",
X"FC18",
X"FC18",
X"FE0C",
X"01F4",
X"0753",
X"0DAC",
X"130B",
X"1388",
X"0E29",
X"02EE",
X"F448",
X"E719",
X"E1BA",
X"E331",
X"E796",
X"ED72",
X"F63C",
X"FF83",
X"0753",
X"0CB2",
X"0F23",
X"0F23",
X"0D2F",
X"0A41",
X"0659",
X"0177",
X"FE0C",
X"FB9B",
X"FB9B",
X"FD8F",
X"0177",
X"06D6",
X"0CB2",
X"128E",
X"1482",
X"0F23",
X"03E8",
X"F542",
X"E813",
X"E237",
X"E3AE",
X"E719",
X"ECF5",
X"F542",
X"FF83",
X"0753",
X"0D2F",
X"0FA0",
X"0F23",
X"0D2F",
X"0A41",
X"05DC",
X"00FA",
X"FD12",
X"FB1E",
X"FB1E",
X"FD8F",
X"00FA",
X"06D6",
X"0D2F",
X"1388",
X"15F9",
X"101D",
X"036B",
X"F34E",
X"E69C",
X"E1BA",
X"E2B4",
X"E69C",
X"ECF5",
X"F63C",
X"0000",
X"084D",
X"0E29",
X"101D",
X"0FA0",
X"0E29",
X"0ABE",
X"055F",
X"007D",
X"FD12",
X"FAA1",
X"FAA1",
X"FC95",
X"00FA",
X"0659",
X"0DAC",
X"1482",
X"16F3",
X"101D",
X"01F4",
X"F15A",
X"E4A8",
X"E0C0",
X"E237",
X"E61F",
X"EDEF",
X"F7B3",
X"0177",
X"09C4",
X"0FA0",
X"1117",
X"109A",
X"0EA6",
X"0ABE",
X"04E2",
X"FF83",
X"FC18",
X"FA24",
X"FA24",
X"FC18",
X"00FA",
X"0659",
X"0DAC",
X"157C",
X"17ED",
X"1117",
X"01F4",
X"F060",
X"E4A8",
X"E043",
X"E1BA",
X"E5A2",
X"ED72",
X"F7B3",
X"01F4",
X"0ABE",
X"101D",
X"1194",
X"109A",
X"0EA6",
X"0ABE",
X"04E2",
X"FF06",
X"FB9B",
X"FA24",
X"FA24",
X"FC95",
X"00FA",
X"0659",
X"0DAC",
X"15F9",
X"186A",
X"1117",
X"007D",
X"EE6C",
X"E3AE",
X"E043",
X"E1BA",
X"E5A2",
X"EE6C",
X"F92A",
X"036B",
X"0BB8",
X"101D",
X"1117",
X"101D",
X"0F23",
X"0ABE",
X"04E2",
X"FF83",
X"FC18",
X"FA24",
X"F92A",
X"FB1E",
X"0000",
X"0659",
X"0DAC",
X"15F9",
X"18E7",
X"1117",
X"0000",
X"ED72",
X"E331",
X"E0C0",
X"E1BA",
X"E5A2",
X"EEE9",
X"FA24",
X"036B",
X"0ABE",
X"0F23",
X"101D",
X"101D",
X"0F23",
X"0BB8",
X"05DC",
X"007D",
X"FC95",
X"FAA1",
X"F8AD",
X"FAA1",
X"0000",
X"06D6",
X"0EA6",
X"16F3",
X"1A5E",
X"1194",
X"FE0C",
X"EB7E",
X"E331",
X"E0C0",
X"E0C0",
X"E5A2",
X"EFE3",
X"FAA1",
X"03E8",
X"0BB8",
X"101D",
X"109A",
X"109A",
X"0F23",
X"0B3B",
X"055F",
X"007D",
X"FC95",
X"F9A7",
X"F830",
X"FAA1",
X"FF83",
X"0659",
X"0FA0",
X"18E7",
X"1ADB",
X"0FA0",
X"FAA1",
X"E90D",
X"E1BA",
X"E043",
X"E043",
X"E69C",
X"F1D7",
X"FC95",
X"055F",
X"0CB2",
X"1117",
X"1194",
X"1117",
X"0EA6",
X"09C4",
X"0465",
X"0000",
X"FC18",
X"F8AD",
X"F736",
X"FAA1",
X"007D",
X"084D",
X"128E",
X"1C52",
X"1C52",
X"0DAC",
X"F6B9",
X"E61F",
X"DFC6",
X"DDD2",
X"DECC",
X"E719",
X"F2D1",
X"FD8F",
X"0753",
X"0FA0",
X"130B",
X"1388",
X"1211",
X"0E29",
X"07D0",
X"01F4",
X"FD8F",
X"FA24",
X"F7B3",
X"F736",
X"FB9B",
X"01F4",
X"0ABE",
X"157C",
X"1FBD",
X"1DC9",
X"0C35",
X"F3CB",
X"E4A8",
X"DFC6",
X"DC5B",
X"DD55",
X"E61F",
X"F34E",
X"FE0C",
X"084D",
X"109A",
X"130B",
X"130B",
X"1194",
X"0E29",
X"07D0",
X"01F4",
X"FD8F",
X"FB1E",
X"F92A",
X"F8AD",
X"FC18",
X"0271",
X"0BB8",
X"1770",
X"203A",
X"1B58",
X"07D0",
X"EFE3",
X"E3AE",
X"DF49",
X"DC5B",
X"DDD2",
X"E813",
X"F542",
X"FF83",
X"09C4",
X"109A",
X"128E",
X"128E",
X"1117",
X"0D2F",
X"06D6",
X"0177",
X"FE0C",
X"FB1E",
X"F8AD",
X"F92A",
X"FC95",
X"0465",
X"0E29",
X"1A5E",
X"20B7",
X"18E7",
X"01F4",
X"EB01",
X"E13D",
X"DD55",
X"DB61",
X"DF49",
X"EBFB",
X"F92A",
X"02EE",
X"0C35",
X"1117",
X"1211",
X"1194",
X"101D",
X"0B3B",
X"055F",
X"007D",
X"FD8F",
X"FA24",
X"F830",
X"F92A",
X"FE89",
X"0753",
X"1194",
X"1DC9",
X"21B1",
X"157C",
X"FB1E",
X"E61F",
X"DF49",
X"DBDE",
X"DA67",
X"E043",
X"EF66",
X"FC18",
X"05DC",
X"0EA6",
X"1211",
X"130B",
X"1211",
X"0F23",
X"09C4",
X"03E8",
X"FF06",
X"FC18",
X"F9A7",
X"F8AD",
X"FAA1",
X"007D",
X"0947",
X"1482",
X"20B7",
X"203A",
X"0F23",
X"F2D1",
X"E2B4",
X"DECC",
X"DAE4",
X"DA67",
X"E42B",
X"F3CB",
X"FF06",
X"09C4",
X"1117",
X"130B",
X"130B",
X"1211",
X"0D2F",
X"0753",
X"0177",
X"FD12",
X"FAA1",
X"F8AD",
X"F92A",
X"FB1E",
X"0177",
X"0B3B",
X"19E1",
X"2422",
X"1E46",
X"07D0",
X"EC78",
X"E1BA",
X"DCD8",
X"D96D",
X"DB61",
X"E90D",
X"F830",
X"0271",
X"0D2F",
X"130B",
X"1388",
X"1388",
X"1194",
X"0BB8",
X"04E2",
X"FE89",
X"FB9B",
X"F9A7",
X"F830",
X"F8AD",
X"FC18",
X"036B",
X"0F23",
X"1EC3",
X"23A5",
X"17ED",
X"FD12",
X"E813",
X"E1BA",
X"DC5B",
X"D96D",
X"DECC",
X"EEE9",
X"FB9B",
X"0659",
X"109A",
X"1405",
X"1482",
X"1405",
X"0FA0",
X"08CA",
X"01F4",
X"FB9B",
X"F9A7",
X"F8AD",
X"F830",
X"F9A7",
X"FD8F",
X"06D6",
X"15F9",
X"23A5",
X"2134",
X"0F23",
X"F2D1",
X"E525",
X"DFC6",
X"DAE4",
X"D9EA",
X"E42B",
X"F448",
X"FF83",
X"0B3B",
X"130B",
X"1388",
X"1482",
X"130B",
X"0DAC",
X"0659",
X"FF06",
X"FA24",
X"FA24",
X"F92A",
X"F8AD",
X"FA24",
X"0000",
X"0B3B",
X"1D4C",
X"2616",
X"1C52",
X"036B",
X"EB01",
X"E3AE",
X"DD55",
X"D7F6",
X"DAE4",
X"EA84",
X"F92A",
X"0465",
X"0FA0",
X"1388",
X"1405",
X"157C",
X"1194",
X"0ABE",
X"02EE",
X"FC18",
X"F9A7",
X"F9A7",
X"F830",
X"F7B3",
X"FAA1",
X"036B",
X"130B",
X"251C",
X"251C",
X"1482",
X"F736",
X"E719",
X"E1BA",
X"DAE4",
X"D873",
X"E043",
X"F0DD",
X"FD12",
X"084D",
X"1194",
X"130B",
X"157C",
X"14FF",
X"0EA6",
X"0753",
X"FF83",
X"FA24",
X"F9A7",
X"F92A",
X"F7B3",
X"F7B3",
X"FE0C",
X"09C4",
X"1DC9",
X"2981",
X"20B7",
X"0753",
X"EBFB",
X"E3AE",
X"DD55",
X"D7F6",
X"D9EA",
X"E890",
X"F7B3",
X"01F4",
X"0E29",
X"1388",
X"1388",
X"15F9",
X"128E",
X"0A41",
X"0271",
X"FB9B",
X"F8AD",
X"F9A7",
X"F92A",
X"F8AD",
X"FAA1",
X"02EE",
X"128E",
X"278D",
X"2904",
X"1676",
X"F7B3",
X"E61F",
X"E13D",
X"D96D",
X"D6FC",
X"DF49",
X"F15A",
X"FE0C",
X"07D0",
X"1211",
X"128E",
X"128E",
X"128E",
X"0D2F",
X"0659",
X"0000",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F9A7",
X"FE0C",
X"0947",
X"1EC3",
X"2CEC",
X"2328",
X"07D0",
X"EB7E",
X"E42B",
X"DD55",
X"D67F",
X"D873",
X"E796",
X"F92A",
X"02EE",
X"0FA0",
X"1482",
X"130B",
X"1388",
X"0F23",
X"08CA",
X"01F4",
X"FB9B",
X"F830",
X"F830",
X"F830",
X"F9A7",
X"FC95",
X"036B",
X"14FF",
X"2AF8",
X"2AF8",
X"1676",
X"F448",
X"E42B",
X"E0C0",
X"D96D",
X"D602",
X"DE4F",
X"F2D1",
X"FF83",
X"0A41",
X"1405",
X"1388",
X"1482",
X"128E",
X"0B3B",
X"04E2",
X"FD8F",
X"F7B3",
X"F5BF",
X"F736",
X"F92A",
X"FB9B",
X"007D",
X"09C4",
X"22AB",
X"2E63",
X"23A5",
X"03E8",
X"E890",
X"E1BA",
X"DB61",
X"D602",
X"D779",
X"EB01",
X"FC95",
X"06D6",
X"1405",
X"15F9",
X"1388",
X"130B",
X"0C35",
X"04E2",
X"FF06",
X"F8AD",
X"F5BF",
X"F830",
X"FA24",
X"FB9B",
X"00FA",
X"04E2",
X"17ED",
X"2C6F",
X"2887",
X"109A",
X"EE6C",
X"E2B4",
X"DCD8",
X"D8F0",
X"D6FC",
X"E525",
X"FB9B",
X"05DC",
X"101D",
X"15F9",
X"128E",
X"1211",
X"0D2F",
X"0465",
X"FF83",
X"FB1E",
X"F6B9",
X"F736",
X"FA24",
X"FC18",
X"0000",
X"0465",
X"0CB2",
X"2599",
X"2A7B",
X"1ADB",
X"F7B3",
X"E331",
X"DECC",
X"DAE4",
X"D9EA",
X"E043",
X"F736",
X"04E2",
X"0CB2",
X"157C",
X"1388",
X"109A",
X"0EA6",
X"06D6",
X"0000",
X"FD12",
X"F8AD",
X"F6B9",
X"F830",
X"FB9B",
X"FE0C",
X"02EE",
X"0659",
X"1BD5",
X"2BF2",
X"222E",
X"055F",
X"E61F",
X"DF49",
X"DB61",
X"DBDE",
X"DC5B",
X"EE6C",
X"0271",
X"09C4",
X"130B",
X"157C",
X"1117",
X"101D",
X"0A41",
X"0177",
X"FD12",
X"F8AD",
X"F5BF",
X"F6B9",
X"FA24",
X"FE89",
X"02EE",
X"05DC",
X"130B",
X"29FE",
X"2693",
X"109A",
X"ECF5",
X"DECC",
X"DB61",
X"DCD8",
X"DD55",
X"E719",
X"FE89",
X"09C4",
X"109A",
X"15F9",
X"1194",
X"0F23",
X"0BB8",
X"03E8",
X"FD12",
X"F92A",
X"F63C",
X"F6B9",
X"F92A",
X"FE89",
X"0271",
X"0753",
X"0C35",
X"23A5",
X"2887",
X"186A",
X"F7B3",
X"DECC",
X"DA67",
X"DB61",
X"DFC6",
X"E331",
X"F830",
X"0947",
X"0EA6",
X"157C",
X"1388",
X"0F23",
X"0C35",
X"05DC",
X"FE89",
X"FAA1",
X"F6B9",
X"F63C",
X"F92A",
X"FE0C",
X"01F4",
X"06D6",
X"0947",
X"1A5E",
X"29FE",
X"1CCF",
X"036B",
X"E2B4",
X"D9EA",
X"D96D",
X"E043",
X"E331",
X"F060",
X"0659",
X"0E29",
X"1388",
X"1676",
X"109A",
X"0CB2",
X"05DC",
X"007D",
X"FB1E",
X"F8AD",
X"F6B9",
X"F7B3",
X"FB9B",
X"007D",
X"055F",
X"08CA",
X"1388",
X"2A7B",
X"222E",
X"0C35",
X"EA84",
X"D8F0",
X"D779",
X"DCD8",
X"E42B",
X"EA07",
X"0177",
X"0E29",
X"1117",
X"15F9",
X"1211",
X"0D2F",
X"0753",
X"0177",
X"FC95",
X"F9A7",
X"F830",
X"F7B3",
X"FA24",
X"FF06",
X"036B",
X"0A41",
X"0EA6",
X"2422",
X"280A",
X"1211",
X"F448",
X"D8F0",
X"D6FC",
X"D9EA",
X"E61F",
X"EA07",
X"F92A",
X"0DAC",
X"1117",
X"1482",
X"128E",
X"0CB2",
X"08CA",
X"02EE",
X"FF06",
X"F9A7",
X"F830",
X"F830",
X"FA24",
X"FD12",
X"007D",
X"084D",
X"0CB2",
X"1BD5",
X"2BF2",
X"18E7",
X"FF83",
X"DECC",
X"D508",
X"D67F",
X"E331",
X"EBFB",
X"F254",
X"09C4",
X"1388",
X"1405",
X"130B",
X"0D2F",
X"09C4",
X"036B",
X"0000",
X"FC95",
X"F7B3",
X"F6B9",
X"F830",
X"FC18",
X"00FA",
X"0753",
X"0CB2",
X"1405",
X"2AF8",
X"20B7",
X"055F",
X"E61F",
X"D391",
X"D585",
X"DE4F",
X"ECF5",
X"F0DD",
X"02EE",
X"1405",
X"1405",
X"130B",
X"0EA6",
X"09C4",
X"0465",
X"FF83",
X"FE0C",
X"F92A",
X"F542",
X"F63C",
X"F9A7",
X"0177",
X"084D",
X"0F23",
X"1194",
X"2599",
X"251C",
X"08CA",
X"ECF5",
X"D40E",
X"D40E",
X"DBDE",
X"EC78",
X"F448",
X"FE0C",
X"1211",
X"157C",
X"128E",
X"0F23",
X"08CA",
X"03E8",
X"FC95",
X"FAA1",
X"F9A7",
X"F6B9",
X"F736",
X"FAA1",
X"0271",
X"0947",
X"0FA0",
X"1117",
X"1DC9",
X"29FE",
X"0EA6",
X"F34E",
X"D779",
X"D120",
X"D873",
X"E813",
X"F5BF",
X"FB9B",
X"0F23",
X"186A",
X"1405",
X"0F23",
X"07D0",
X"036B",
X"FE89",
X"FAA1",
X"F92A",
X"F736",
X"F830",
X"FC95",
X"007D",
X"06D6",
X"0C35",
X"0EA6",
X"157C",
X"2AF8",
X"1B58",
X"FC18",
X"E0C0",
X"CFA9",
X"D40E",
X"E0C0",
X"F2D1",
X"F92A",
X"0947",
X"1A5E",
X"18E7",
X"1117",
X"07D0",
X"0177",
X"FE0C",
X"F92A",
X"F8AD",
X"F92A",
X"F830",
X"FE89",
X"00FA",
X"036B",
X"0947",
X"0EA6",
X"1117",
X"2616",
X"251C",
X"036B",
X"E890",
X"D026",
X"D0A3",
X"DBDE",
X"EEE9",
X"F9A7",
X"03E8",
X"1770",
X"1BD5",
X"157C",
X"0ABE",
X"02EE",
X"FF06",
X"FA24",
X"F736",
X"F8AD",
X"F830",
X"FB9B",
X"007D",
X"0271",
X"07D0",
X"0E29",
X"0F23",
X"1DC9",
X"2A7B",
X"0ABE",
X"EEE9",
X"D602",
X"CEAF",
X"D8F0",
X"EA07",
X"FA24",
X"FF83",
X"0F23",
X"1964",
X"186A",
X"0EA6",
X"03E8",
X"00FA",
X"FC95",
X"F8AD",
X"FA24",
X"FB9B",
X"FB1E",
X"FF06",
X"007D",
X"0271",
X"0A41",
X"0EA6",
X"14FF",
X"2BF2",
X"17ED",
X"F5BF",
X"DECC",
X"CF2C",
X"D67F",
X"E3AE",
X"F736",
X"FD8F",
X"084D",
X"16F3",
X"18E7",
X"128E",
X"036B",
X"FF83",
X"FF06",
X"FB9B",
X"FC95",
X"0000",
X"FE0C",
X"FE89",
X"FE0C",
X"FF06",
X"04E2",
X"0CB2",
X"0C35",
X"251C",
X"2710",
X"007D",
X"E890",
X"D297",
X"D297",
X"DECC",
X"F1D7",
X"FE89",
X"01F4",
X"1117",
X"17ED",
X"1405",
X"0753",
X"FE89",
X"00FA",
X"FE89",
X"FAA1",
X"FD12",
X"FE0C",
X"0000",
X"0000",
X"FF06",
X"01F4",
X"0BB8",
X"0BB8",
X"1676",
X"2DE6",
X"0F23",
X"EEE9",
X"D96D",
X"D19D",
X"DBDE",
X"EB01",
X"FD8F",
X"007D",
X"09C4",
X"186A",
X"17ED",
X"0CB2",
X"FF83",
X"00FA",
X"007D",
X"F8AD",
X"F7B3",
X"F8AD",
X"FC95",
X"0465",
X"00FA",
X"00FA",
X"0A41",
X"101D",
X"0C35",
X"278D",
X"1F40",
X"F63C",
X"DECC",
X"D026",
X"D67F",
X"E4A8",
X"FA24",
X"036B",
X"0465",
X"130B",
X"18E7",
X"109A",
X"02EE",
X"FE0C",
X"02EE",
X"FC18",
X"F7B3",
X"F830",
X"FA24",
X"00FA",
X"036B",
X"0271",
X"0753",
X"1405",
X"0E29",
X"18E7",
X"278D",
X"036B",
X"E61F",
X"D391",
X"D21A",
X"DD55",
X"F3CB",
X"04E2",
X"036B",
X"0CB2",
X"186A",
X"1388",
X"06D6",
X"FB9B",
X"00FA",
X"0000",
X"F92A",
X"F830",
X"F8AD",
X"FC95",
X"01F4",
X"04E2",
X"05DC",
X"109A",
X"14FF",
X"0D2F",
X"2422",
X"15F9",
X"F254",
X"DAE4",
X"D19D",
X"D6FC",
X"E719",
X"FF83",
X"036B",
X"04E2",
X"15F9",
X"1770",
X"101D",
X"01F4",
X"FC95",
X"007D",
X"FB9B",
X"F830",
X"F736",
X"FA24",
X"FE89",
X"01F4",
X"0659",
X"0BB8",
X"186A",
X"0D2F",
X"1676",
X"222E",
X"036B",
X"E719",
X"D48B",
X"D48B",
X"DCD8",
X"F4C5",
X"04E2",
X"0177",
X"0CB2",
X"1770",
X"1388",
X"0947",
X"FC95",
X"007D",
X"0000",
X"FB1E",
X"F830",
X"F92A",
X"FB9B",
X"00FA",
X"03E8",
X"0659",
X"109A",
X"1211",
X"09C4",
X"21B1",
X"1770",
X"F542",
X"DCD8",
X"D508",
X"D779",
X"E719",
X"FF83",
X"04E2",
X"055F",
X"14FF",
X"16F3",
X"0F23",
X"01F4",
X"FC18",
X"00FA",
X"FE0C",
X"F92A",
X"F9A7",
X"FA24",
X"00FA",
X"0465",
X"01F4",
X"0659",
X"1117",
X"084D",
X"128E",
X"251C",
X"09C4",
X"EA07",
X"D8F0",
X"D779",
X"DC5B",
X"F3CB",
X"03E8",
X"036B",
X"0D2F",
X"186A",
X"1388",
X"09C4",
X"FC18",
X"FD8F",
X"007D",
X"FB9B",
X"F9A7",
X"F9A7",
X"FB9B",
X"02EE",
X"01F4",
X"007D",
X"09C4",
X"0EA6",
X"0753",
X"1F40",
X"1B58",
X"FA24",
X"DECC",
X"D6FC",
X"DA67",
X"E890",
X"00FA",
X"084D",
X"084D",
X"130B",
X"1405",
X"0DAC",
X"FF83",
X"F830",
X"FF06",
X"FE0C",
X"FB1E",
X"FD12",
X"FF83",
X"0000",
X"0177",
X"0177",
X"007D",
X"09C4",
X"05DC",
X"0F23",
X"22AB",
X"0E29",
X"F1D7",
X"DA67",
X"DA67",
X"E0C0",
X"F3CB",
X"06D6",
X"06D6",
X"0BB8",
X"128E",
X"0EA6",
X"07D0",
X"FB1E",
X"FB1E",
X"FE89",
X"FB9B",
X"F92A",
X"FB1E",
X"FE89",
X"0177",
X"036B",
X"0177",
X"06D6",
X"0D2F",
X"05DC",
X"18E7",
X"1BD5",
X"036B",
X"E90D",
X"D873",
X"DDD2",
X"EA07",
X"FE89",
X"0947",
X"07D0",
X"0FA0",
X"128E",
X"0C35",
X"0271",
X"F92A",
X"FC18",
X"FB9B",
X"FA24",
X"F8AD",
X"FB9B",
X"00FA",
X"03E8",
X"0271",
X"0271",
X"0947",
X"0947",
X"09C4",
X"1C52",
X"1388",
X"FB1E",
X"E237",
X"D9EA",
X"E42B",
X"F254",
X"0271",
X"05DC",
X"04E2",
X"101D",
X"0FA0",
X"0ABE",
X"FF83",
X"F92A",
X"FD8F",
X"FC95",
X"FC95",
X"FC95",
X"FE0C",
X"01F4",
X"02EE",
X"007D",
X"0271",
X"07D0",
X"05DC",
X"0E29",
X"1D4C",
X"0F23",
X"F3CB",
X"DDD2",
X"DF49",
X"E98A",
X"F7B3",
X"0465",
X"0465",
X"06D6",
X"0F23",
X"0ABE",
X"0659",
X"FD8F",
X"FB1E",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE89",
X"01F4",
X"0177",
X"0000",
X"036B",
X"07D0",
X"0659",
X"130B",
X"1B58",
X"08CA",
X"EC78",
X"DD55",
X"E13D",
X"EA84",
X"F9A7",
X"036B",
X"0465",
X"0BB8",
X"101D",
X"0BB8",
X"05DC",
X"FC95",
X"FC18",
X"FE0C",
X"FE89",
X"FD12",
X"FD8F",
X"0000",
X"02EE",
X"007D",
X"00FA",
X"06D6",
X"07D0",
X"08CA",
X"16F3",
X"18E7",
X"055F",
X"EA07",
X"DE4F",
X"E13D",
X"EC78",
X"FB9B",
X"0177",
X"0465",
X"0CB2",
X"0EA6",
X"0ABE",
X"036B",
X"FC18",
X"FD12",
X"FF06",
X"FD8F",
X"FB1E",
X"FE0C",
X"0000",
X"FF83",
X"FE89",
X"00FA",
X"0659",
X"07D0",
X"0BB8",
X"1770",
X"157C",
X"FF83",
X"E796",
X"E043",
X"E525",
X"F0DD",
X"FD8F",
X"02EE",
X"0753",
X"0D2F",
X"0CB2",
X"0947",
X"01F4",
X"FD12",
X"FE89",
X"FE89",
X"FB9B",
X"FA24",
X"FB9B",
X"FD8F",
X"00FA",
X"01F4",
X"04E2",
X"0A41",
X"0A41",
X"0F23",
X"17ED",
X"0F23",
X"F9A7",
X"E719",
X"E2B4",
X"E719",
X"F1D7",
X"FD12",
X"007D",
X"05DC",
X"0A41",
X"0B3B",
X"07D0",
X"00FA",
X"FE0C",
X"FE89",
X"FF06",
X"FC18",
X"FC18",
X"FD8F",
X"FF83",
X"0177",
X"0271",
X"06D6",
X"0ABE",
X"0ABE",
X"1194",
X"1482",
X"084D",
X"F542",
X"E719",
X"E4A8",
X"E98A",
X"F63C",
X"FF06",
X"036B",
X"084D",
X"0A41",
X"0B3B",
X"0753",
X"007D",
X"FD8F",
X"FE0C",
X"FE0C",
X"FB9B",
X"FC18",
X"FD8F",
X"FF06",
X"007D",
X"036B",
X"06D6",
X"09C4",
X"0B3B",
X"130B",
X"1211",
X"05DC",
X"F4C5",
X"E90D",
X"E525",
X"EA07",
X"F63C",
X"FD8F",
X"03E8",
X"06D6",
X"084D",
X"0947",
X"05DC",
X"0177",
X"FF06",
X"FE89",
X"FF06",
X"FD12",
X"FD12",
X"FD8F",
X"FF83",
X"007D",
X"036B",
X"0753",
X"09C4",
X"0CB2",
X"130B",
X"0E29",
X"01F4",
X"F4C5",
X"EB7E",
X"E813",
X"ED72",
X"F5BF",
X"FE89",
X"0659",
X"084D",
X"08CA",
X"06D6",
X"036B",
X"0000",
X"FF06",
X"FF06",
X"FE0C",
X"FD8F",
X"FD12",
X"FE89",
X"007D",
X"007D",
X"02EE",
X"0659",
X"0947",
X"0DAC",
X"128E",
X"0B3B",
X"007D",
X"F542",
X"ECF5",
X"EA84",
X"EE6C",
X"F542",
X"FE0C",
X"04E2",
X"084D",
X"08CA",
X"0753",
X"02EE",
X"0000",
X"FF06",
X"FE0C",
X"FE0C",
X"FD8F",
X"FE89",
X"007D",
X"00FA",
X"007D",
X"0271",
X"055F",
X"0753",
X"0ABE",
X"0B3B",
X"0465",
X"FF83",
X"F8AD",
X"F3CB",
X"F254",
X"F254",
X"F542",
X"FB1E",
X"007D",
X"0465",
X"0753",
X"0753",
X"04E2",
X"03E8",
X"01F4",
X"007D",
X"FF83",
X"FE0C",
X"FE89",
X"0000",
X"007D",
X"00FA",
X"02EE",
X"04E2",
X"05DC",
X"07D0",
X"055F",
X"0000",
X"FC18",
X"F830",
X"F7B3",
X"F92A",
X"F92A",
X"F92A",
X"FB9B",
X"FE0C",
X"00FA",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"02EE",
X"0177",
X"FF83",
X"FE0C",
X"FE0C",
X"FF83",
X"0000",
X"00FA",
X"036B",
X"055F",
X"06D6",
X"0753",
X"03E8",
X"0000",
X"FC18",
X"F92A",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FC18",
X"FE0C",
X"007D",
X"0271",
X"036B",
X"03E8",
X"03E8",
X"02EE",
X"0177",
X"FF06",
X"FE0C",
X"FE0C",
X"FF06",
X"FF83",
X"00FA",
X"036B",
X"055F",
X"0753",
X"0659",
X"02EE",
X"0000",
X"FB9B",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"FAA1",
X"FC18",
X"FE0C",
X"00FA",
X"0271",
X"03E8",
X"04E2",
X"04E2",
X"036B",
X"00FA",
X"FE89",
X"FD12",
X"FE0C",
X"FE89",
X"FF06",
X"007D",
X"02EE",
X"05DC",
X"07D0",
X"05DC",
X"0271",
X"FF83",
X"FC95",
X"FB9B",
X"FB1E",
X"FA24",
X"F9A7",
X"FA24",
X"FB9B",
X"FE89",
X"00FA",
X"0271",
X"0465",
X"055F",
X"055F",
X"03E8",
X"00FA",
X"FE0C",
X"FD12",
X"FD12",
X"FD8F",
X"FF06",
X"00FA",
X"03E8",
X"06D6",
X"06D6",
X"03E8",
X"0177",
X"FE89",
X"FC95",
X"FB1E",
X"FA24",
X"F92A",
X"FA24",
X"FB9B",
X"FD12",
X"FF06",
X"00FA",
X"0271",
X"03E8",
X"04E2",
X"0465",
X"036B",
X"0177",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FF83",
X"007D",
X"02EE",
X"04E2",
X"0465",
X"01F4",
X"007D",
X"FE89",
X"FD8F",
X"FC18",
X"FB1E",
X"FAA1",
X"FB9B",
X"FC95",
X"FE89",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"02EE",
X"0271",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FF83",
X"0000",
X"0177",
X"036B",
X"04E2",
X"036B",
X"0177",
X"FF83",
X"FE0C",
X"FD8F",
X"FC95",
X"FB9B",
X"FB9B",
X"FC18",
X"FD12",
X"FE0C",
X"FF83",
X"007D",
X"0177",
X"02EE",
X"036B",
X"02EE",
X"0271",
X"0177",
X"007D",
X"FF83",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"02EE",
X"036B",
X"0271",
X"00FA",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"0177",
X"02EE",
X"02EE",
X"02EE",
X"01F4",
X"0177",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"0177",
X"02EE",
X"02EE",
X"0271",
X"00FA",
X"FF83",
X"FE89",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FF83",
X"0177",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"007D",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"00FA",
X"01F4",
X"0271",
X"01F4",
X"00FA",
X"0000",
X"FE89",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"007D",
X"01F4",
X"036B",
X"02EE",
X"0271",
X"0271",
X"0177",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"0177",
X"0177",
X"0177",
X"007D",
X"FF83",
X"FE0C",
X"FD8F",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FF06",
X"0000",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"0177",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FD8F",
X"FD12",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF83",
X"007D",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"0000",
X"007D",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"01F4",
X"0271",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"01F4",
X"01F4",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"01F4",
X"0271",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE89",
X"FF83",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"00FA",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"0177",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FD8F",
X"FE0C",
X"FF83",
X"007D",
X"0177",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"01F4",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"00FA",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"007D",
X"0177",
X"0271",
X"02EE",
X"036B",
X"02EE",
X"0271",
X"0177",
X"007D",
X"0000",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"0177",
X"007D",
X"0000",
X"FF06",
X"FE0C",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FD8F",
X"FE89",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"036B",
X"02EE",
X"01F4",
X"00FA",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"007D",
X"0177",
X"0271",
X"036B",
X"036B",
X"036B",
X"0271",
X"0177",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FE0C",
X"FF83",
X"00FA",
X"01F4",
X"02EE",
X"03E8",
X"03E8",
X"036B",
X"0271",
X"00FA",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"0000",
X"FE89",
X"FD8F",
X"FD12",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FD8F",
X"FE89",
X"0000",
X"0177",
X"0271",
X"036B",
X"03E8",
X"036B",
X"02EE",
X"01F4",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"0177",
X"01F4",
X"01F4",
X"0177",
X"007D",
X"FF83",
X"FE0C",
X"FD12",
X"FC95",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FE0C",
X"FF83",
X"007D",
X"01F4",
X"02EE",
X"036B",
X"03E8",
X"036B",
X"0271",
X"0177",
X"007D",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD12",
X"FC18",
X"FB9B",
X"FB9B",
X"FC18",
X"FD12",
X"FE89",
X"0000",
X"0177",
X"0271",
X"036B",
X"03E8",
X"03E8",
X"02EE",
X"01F4",
X"00FA",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"00FA",
X"FF83",
X"FE89",
X"FD8F",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FD8F",
X"FF06",
X"007D",
X"01F4",
X"036B",
X"03E8",
X"0465",
X"03E8",
X"02EE",
X"0177",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0177",
X"007D",
X"FF83",
X"FE0C",
X"FD12",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC95",
X"FE0C",
X"FF83",
X"00FA",
X"0271",
X"03E8",
X"0465",
X"0465",
X"036B",
X"0271",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"01F4",
X"0271",
X"0271",
X"0177",
X"007D",
X"FF06",
X"FD8F",
X"FC95",
X"FB9B",
X"FB1E",
X"FB1E",
X"FB9B",
X"FD12",
X"FE89",
X"0000",
X"01F4",
X"02EE",
X"03E8",
X"0465",
X"0465",
X"036B",
X"01F4",
X"007D",
X"FF83",
X"FE89",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"0271",
X"0271",
X"01F4",
X"00FA",
X"FF83",
X"FE89",
X"FD12",
X"FC18",
X"FB1E",
X"FB1E",
X"FB1E",
X"FC18",
X"FD12",
X"FF06",
X"00FA",
X"0271",
X"03E8",
X"0465",
X"04E2",
X"03E8",
X"02EE",
X"0177",
X"0000",
X"FF06",
X"FE89",
X"FF06",
X"FF83",
X"00FA",
X"01F4",
X"0271",
X"0271",
X"01F4",
X"007D",
X"FF06",
X"FD8F",
X"FC95",
X"FB9B",
X"FB1E",
X"FB1E",
X"FB9B",
X"FC95",
X"FE0C",
X"0000",
X"0177",
X"02EE",
X"0465",
X"04E2",
X"04E2",
X"03E8",
X"0271",
X"00FA",
X"FF83",
X"FF06",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"01F4",
X"0271",
X"0271",
X"0177",
X"0000",
X"FE89",
X"FD12",
X"FC18",
X"FB1E",
X"FAA1",
X"FB1E",
X"FB9B",
X"FD12",
X"FE89",
X"007D",
X"0271",
X"03E8",
X"04E2",
X"04E2",
X"0465",
X"036B",
X"01F4",
X"007D",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"007D",
X"0177",
X"0271",
X"0271",
X"01F4",
X"00FA",
X"FF83",
X"FE0C",
X"FC95",
X"FB9B",
X"FAA1",
X"FAA1",
X"FB1E",
X"FC18",
X"FD8F",
X"FF83",
X"0177",
X"02EE",
X"0465",
X"055F",
X"055F",
X"0465",
X"02EE",
X"0177",
X"0000",
X"FE89",
X"FE0C",
X"FE89",
X"FF83",
X"007D",
X"01F4",
X"02EE",
X"0271",
X"01F4",
X"007D",
X"FF06",
X"FD8F",
X"FC18",
X"FB1E",
X"FAA1",
X"FAA1",
X"FAA1",
X"FC18",
X"FD8F",
X"0000",
X"01F4",
X"036B",
X"04E2",
X"055F",
X"055F",
X"0465",
X"02EE",
X"00FA",
X"FF83",
X"FE89",
X"FE0C",
X"FE89",
X"0000",
X"00FA",
X"0271",
X"02EE",
X"02EE",
X"01F4",
X"0000",
X"FE89",
X"FD12",
X"FB9B",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FC18",
X"FE89",
X"007D",
X"0271",
X"0465",
X"055F",
X"05DC",
X"055F",
X"0465",
X"0271",
X"007D",
X"FF06",
X"FE0C",
X"FE0C",
X"FE89",
X"0000",
X"01F4",
X"02EE",
X"036B",
X"02EE",
X"0177",
X"FF83",
X"FE0C",
X"FC95",
X"FB1E",
X"FA24",
X"F9A7",
X"FA24",
X"FB1E",
X"FC95",
X"FF06",
X"00FA",
X"036B",
X"04E2",
X"05DC",
X"05DC",
X"055F",
X"03E8",
X"01F4",
X"0000",
X"FE89",
X"FD8F",
X"FE0C",
X"FF06",
X"00FA",
X"0271",
X"036B",
X"036B",
X"02EE",
X"00FA",
X"FF06",
X"FD8F",
X"FC18",
X"FAA1",
X"F9A7",
X"F9A7",
X"F9A7",
X"FB1E",
X"FD12",
X"FF83",
X"01F4",
X"03E8",
X"055F",
X"0659",
X"05DC",
X"04E2",
X"036B",
X"0177",
X"FF83",
X"FE0C",
X"FD8F",
X"FE0C",
X"FF83",
X"0177",
X"02EE",
X"03E8",
X"03E8",
X"0271",
X"007D",
X"FE89",
X"FD12",
X"FB1E",
X"F9A7",
X"F92A",
X"F92A",
X"F9A7",
X"FB9B",
X"FE0C",
X"007D",
X"0271",
X"0465",
X"05DC",
X"0659",
X"05DC",
X"0465",
X"0271",
X"007D",
X"FF06",
X"FE0C",
X"FD8F",
X"FE89",
X"0000",
X"01F4",
X"036B",
X"0465",
X"03E8",
X"01F4",
X"0000",
X"FE0C",
X"FC95",
X"FAA1",
X"F92A",
X"F92A",
X"F92A",
X"FA24",
X"FC18",
X"FE89",
X"00FA",
X"036B",
X"04E2",
X"0659",
X"0659",
X"055F",
X"03E8",
X"01F4",
X"0000",
X"FE89",
X"FE0C",
X"FE0C",
X"FE89",
X"007D",
X"0271",
X"03E8",
X"0465",
X"036B",
X"0177",
X"FF83",
X"FD8F",
X"FB9B",
X"FA24",
X"F92A",
X"F92A",
X"F9A7",
X"FB1E",
X"FD12",
X"FF83",
X"0177",
X"03E8",
X"055F",
X"0659",
X"0659",
X"055F",
X"036B",
X"0177",
X"FF83",
X"FE0C",
X"FD8F",
X"FD8F",
X"FF06",
X"00FA",
X"02EE",
X"0465",
X"0465",
X"02EE",
X"007D",
X"FE89",
X"FD12",
X"FB1E",
X"F9A7",
X"F92A",
X"F92A",
X"F9A7",
X"FB9B",
X"FD8F",
X"0000",
X"0271",
X"0465",
X"05DC",
X"0659",
X"05DC",
X"04E2",
X"02EE",
X"00FA",
X"FF06",
X"FE0C",
X"FD8F",
X"FE0C",
X"FF83",
X"01F4",
X"03E8",
X"04E2",
X"03E8",
X"01F4",
X"0000",
X"FE0C",
X"FC18",
X"FAA1",
X"F92A",
X"F8AD",
X"F92A",
X"FA24",
X"FC18",
X"FE89",
X"00FA",
X"036B",
X"055F",
X"0659",
X"0659",
X"05DC",
X"0465",
X"0271",
X"007D",
X"FE89",
X"FD8F",
X"FD8F",
X"FE0C",
X"0000",
X"0271",
X"0465",
X"04E2",
X"036B",
X"00FA",
X"FF83",
X"FD8F",
X"FB9B",
X"F9A7",
X"F8AD",
X"F8AD",
X"F92A",
X"FAA1",
X"FD12",
X"FF83",
X"01F4",
X"03E8",
X"05DC",
X"0659",
X"0659",
X"055F",
X"03E8",
X"01F4",
X"0000",
X"FE0C",
X"FD8F",
X"FD8F",
X"FE89",
X"00FA",
X"036B",
X"04E2",
X"0465",
X"0271",
X"007D",
X"FF06",
X"FD12",
X"FB1E",
X"F92A",
X"F8AD",
X"F830",
X"F92A",
X"FB1E",
X"FD8F",
X"0000",
X"0271",
X"04E2",
X"05DC",
X"0659",
X"0659",
X"055F",
X"036B",
X"00FA",
X"FF83",
X"FE0C",
X"FD12",
X"FD8F",
X"FF06",
X"01F4",
X"03E8",
X"04E2",
X"03E8",
X"01F4",
X"0000",
X"FE89",
X"FC95",
X"FA24",
X"F92A",
X"F830",
X"F830",
X"F9A7",
X"FB9B",
X"FE89",
X"00FA",
X"036B",
X"055F",
X"06D6",
X"06D6",
X"0659",
X"04E2",
X"02EE",
X"007D",
X"FE89",
X"FD8F",
X"FD12",
X"FE0C",
X"0000",
X"0271",
X"04E2",
X"04E2",
X"036B",
X"0177",
X"0000",
X"FE0C",
X"FB9B",
X"F9A7",
X"F830",
X"F7B3",
X"F830",
X"FA24",
X"FC95",
X"FF06",
X"01F4",
X"0465",
X"0659",
X"06D6",
X"06D6",
X"0659",
X"0465",
X"01F4",
X"0000",
X"FE0C",
X"FD12",
X"FD12",
X"FE0C",
X"007D",
X"036B",
X"055F",
X"0465",
X"02EE",
X"0177",
X"FF83",
X"FD12",
X"FAA1",
X"F92A",
X"F830",
X"F7B3",
X"F830",
X"FAA1",
X"FD12",
X"0000",
X"02EE",
X"055F",
X"06D6",
X"0753",
X"06D6",
X"05DC",
X"03E8",
X"0177",
X"FF83",
X"FD8F",
X"FD12",
X"FD12",
X"FE89",
X"0177",
X"0465",
X"055F",
X"0465",
X"02EE",
X"0177",
X"FF06",
X"FC18",
X"FA24",
X"F830",
X"F736",
X"F736",
X"F8AD",
X"FB1E",
X"FE0C",
X"007D",
X"036B",
X"05DC",
X"0753",
X"07D0",
X"0753",
X"05DC",
X"036B",
X"00FA",
X"FE89",
X"FD12",
X"FC95",
X"FC95",
X"FF06",
X"01F4",
X"04E2",
X"05DC",
X"0465",
X"02EE",
X"00FA",
X"FE89",
X"FB9B",
X"F92A",
X"F7B3",
X"F6B9",
X"F736",
X"F8AD",
X"FB9B",
X"FE89",
X"0177",
X"0465",
X"06D6",
X"07D0",
X"07D0",
X"06D6",
X"055F",
X"0271",
X"0000",
X"FE0C",
X"FC95",
X"FC18",
X"FD12",
X"FF83",
X"036B",
X"05DC",
X"05DC",
X"0465",
X"0271",
X"007D",
X"FD8F",
X"FAA1",
X"F8AD",
X"F736",
X"F6B9",
X"F7B3",
X"F9A7",
X"FC95",
X"FF83",
X"0271",
X"055F",
X"0753",
X"07D0",
X"07D0",
X"06D6",
X"04E2",
X"01F4",
X"FF83",
X"FD8F",
X"FC18",
X"FC18",
X"FD8F",
X"007D",
X"03E8",
X"05DC",
X"05DC",
X"03E8",
X"01F4",
X"FF83",
X"FC95",
X"FA24",
X"F830",
X"F6B9",
X"F6B9",
X"F7B3",
X"FA24",
X"FD12",
X"0000",
X"036B",
X"05DC",
X"0753",
X"084D",
X"07D0",
X"0659",
X"03E8",
X"00FA",
X"FE89",
X"FC95",
X"FB9B",
X"FC18",
X"FE0C",
X"0177",
X"04E2",
X"0659",
X"05DC",
X"03E8",
X"01F4",
X"FF06",
X"FC18",
X"F9A7",
X"F7B3",
X"F63C",
X"F63C",
X"F7B3",
X"FAA1",
X"FD8F",
X"00FA",
X"03E8",
X"0659",
X"084D",
X"084D",
X"07D0",
X"05DC",
X"036B",
X"007D",
X"FE0C",
X"FC95",
X"FB9B",
X"FC18",
X"FE89",
X"0271",
X"055F",
X"06D6",
X"05DC",
X"03E8",
X"0177",
X"FE89",
X"FB9B",
X"F8AD",
X"F6B9",
X"F5BF",
X"F63C",
X"F830",
X"FB1E",
X"FE0C",
X"0177",
X"04E2",
X"0753",
X"084D",
X"08CA",
X"0753",
X"055F",
X"0271",
X"FF83",
X"FD12",
X"FB9B",
X"FB1E",
X"FC95",
X"FF83",
X"036B",
X"0659",
X"0753",
X"0659",
X"03E8",
X"00FA",
X"FD8F",
X"FAA1",
X"F7B3",
X"F5BF",
X"F542",
X"F63C",
X"F8AD",
X"FB9B",
X"FF06",
X"0271",
X"05DC",
X"084D",
X"0947",
X"08CA",
X"0753",
X"04E2",
X"0177",
X"FE89",
X"FC95",
X"FB1E",
X"FB1E",
X"FD12",
X"007D",
X"0465",
X"0753",
X"07D0",
X"0659",
X"036B",
X"0000",
X"FD12",
X"F92A",
X"F63C",
X"F4C5",
X"F4C5",
X"F63C",
X"F92A",
X"FC95",
X"0000",
X"036B",
X"06D6",
X"08CA",
X"09C4",
X"08CA",
X"06D6",
X"03E8",
X"00FA",
X"FE0C",
X"FB9B",
X"FAA1",
X"FB1E",
X"FD8F",
X"0177",
X"05DC",
X"08CA",
X"084D",
X"05DC",
X"0271",
X"FF06",
X"FB9B",
X"F7B3",
X"F542",
X"F448",
X"F4C5",
X"F6B9",
X"F9A7",
X"FD8F",
X"0177",
X"04E2",
X"084D",
X"09C4",
X"0A41",
X"08CA",
X"06D6",
X"036B",
X"0000",
X"FD12",
X"FAA1",
X"FA24",
X"FB1E",
X"FE0C",
X"01F4",
X"06D6",
X"09C4",
X"08CA",
X"04E2",
X"00FA",
X"FE0C",
X"FAA1",
X"F6B9",
X"F4C5",
X"F448",
X"F4C5",
X"F736",
X"FB1E",
X"FE89",
X"0271",
X"05DC",
X"08CA",
X"0A41",
X"09C4",
X"084D",
X"05DC",
X"02EE",
X"FF06",
X"FC95",
X"FAA1",
X"FA24",
X"FB9B",
X"FE89",
X"036B",
X"07D0",
X"09C4",
X"07D0",
X"03E8",
X"0000",
X"FD12",
X"F92A",
X"F5BF",
X"F448",
X"F448",
X"F542",
X"F830",
X"FB9B",
X"FF83",
X"02EE",
X"06D6",
X"0947",
X"0A41",
X"09C4",
X"07D0",
X"055F",
X"0177",
X"FE0C",
X"FB9B",
X"FA24",
X"FA24",
X"FC18",
X"FF83",
X"04E2",
X"0947",
X"0A41",
X"0753",
X"0271",
X"FF83",
X"FC18",
X"F7B3",
X"F4C5",
X"F3CB",
X"F448",
X"F5BF",
X"F92A",
X"FD12",
X"00FA",
X"04E2",
X"084D",
X"0A41",
X"0A41",
X"0947",
X"0753",
X"0465",
X"0000",
X"FD12",
X"FB1E",
X"FA24",
X"FAA1",
X"FD12",
X"00FA",
X"06D6",
X"0B3B",
X"0ABE",
X"05DC",
X"00FA",
X"FE0C",
X"FAA1",
X"F5BF",
X"F34E",
X"F3CB",
X"F4C5",
X"F6B9",
X"FA24",
X"FE89",
X"0271",
X"05DC",
X"0947",
X"0ABE",
X"0A41",
X"08CA",
X"06D6",
X"02EE",
X"FF06",
X"FC18",
X"FAA1",
X"FA24",
X"FB1E",
X"FE0C",
X"02EE",
X"0947",
X"0C35",
X"09C4",
X"036B",
X"FF83",
X"FD8F",
X"F92A",
X"F3CB",
X"F2D1",
X"F3CB",
X"F448",
X"F736",
X"FB9B",
X"0000",
X"036B",
X"0753",
X"0A41",
X"0ABE",
X"09C4",
X"084D",
X"05DC",
X"0177",
X"FE0C",
X"FB9B",
X"FA24",
X"FA24",
X"FB9B",
X"FF06",
X"04E2",
X"0BB8",
X"0D2F",
X"08CA",
X"0177",
X"FE89",
X"FC18",
X"F63C",
X"F254",
X"F2D1",
X"F3CB",
X"F4C5",
X"F8AD",
X"FD12",
X"0177",
X"04E2",
X"08CA",
X"0ABE",
X"0ABE",
X"0947",
X"0753",
X"03E8",
X"0000",
X"FD12",
X"FAA1",
X"F9A7",
X"FAA1",
X"FD12",
X"00FA",
X"07D0",
X"0DAC",
X"0D2F",
X"05DC",
X"FF06",
X"FE0C",
X"FA24",
X"F3CB",
X"F15A",
X"F3CB",
X"F3CB",
X"F5BF",
X"FAA1",
X"FF83",
X"036B",
X"0659",
X"0A41",
X"0B3B",
X"0A41",
X"08CA",
X"0659",
X"0271",
X"FE89",
X"FB9B",
X"FA24",
X"F9A7",
X"FB1E",
X"FE0C",
X"02EE",
X"0ABE",
X"0EA6",
X"0BB8",
X"0271",
X"FE0C",
X"FD12",
X"F7B3",
X"F1D7",
X"F1D7",
X"F3CB",
X"F448",
X"F736",
X"FC95",
X"00FA",
X"0465",
X"084D",
X"0B3B",
X"0B3B",
X"09C4",
X"08CA",
X"055F",
X"00FA",
X"FD8F",
X"FB9B",
X"F9A7",
X"F92A",
X"FB9B",
X"FE89",
X"0465",
X"0CB2",
X"0FA0",
X"09C4",
X"0000",
X"FE0C",
X"FC18",
X"F4C5",
X"EFE3",
X"F254",
X"F3CB",
X"F3CB",
X"F8AD",
X"FE89",
X"02EE",
X"0659",
X"0A41",
X"0C35",
X"0ABE",
X"0947",
X"0753",
X"036B",
X"FF83",
X"FC95",
X"FAA1",
X"F92A",
X"F9A7",
X"FC95",
X"0000",
X"084D",
X"0FA0",
X"0F23",
X"055F",
X"FD8F",
X"FE0C",
X"F9A7",
X"F1D7",
X"F060",
X"F3CB",
X"F2D1",
X"F4C5",
X"FB9B",
X"00FA",
X"0465",
X"084D",
X"0C35",
X"0BB8",
X"0A41",
X"08CA",
X"05DC",
X"0177",
X"FD8F",
X"FB1E",
X"F9A7",
X"F830",
X"FB1E",
X"FE0C",
X"0271",
X"0D2F",
X"1211",
X"0CB2",
X"FF83",
X"FD12",
X"FE0C",
X"F5BF",
X"EEE9",
X"F1D7",
X"F448",
X"F2D1",
X"F7B3",
X"FF06",
X"02EE",
X"05DC",
X"0A41",
X"0D2F",
X"0B3B",
X"0A41",
X"07D0",
X"03E8",
X"FF83",
X"FB9B",
X"F9A7",
X"F830",
X"F92A",
X"FC95",
X"FE89",
X"07D0",
X"1194",
X"1194",
X"055F",
X"FB9B",
X"FE89",
X"FAA1",
X"F0DD",
X"EEE9",
X"F448",
X"F3CB",
X"F4C5",
X"FC18",
X"0177",
X"0465",
X"0947",
X"0D2F",
X"0C35",
X"09C4",
X"084D",
X"055F",
X"007D",
X"FC95",
X"FAA1",
X"F830",
X"F736",
X"FB1E",
X"FE89",
X"0271",
X"0EA6",
X"1482",
X"0E29",
X"FE89",
X"FB9B",
X"FE0C",
X"F4C5",
X"EC78",
X"F0DD",
X"F542",
X"F2D1",
X"F7B3",
X"0000",
X"03E8",
X"0753",
X"0CB2",
X"0E29",
X"0B3B",
X"0947",
X"06D6",
X"0271",
X"FE0C",
X"FB1E",
X"F830",
X"F63C",
X"F830",
X"FD12",
X"FF06",
X"08CA",
X"1388",
X"130B",
X"0659",
X"FAA1",
X"FE0C",
X"FA24",
X"EF66",
X"ED72",
X"F448",
X"F3CB",
X"F448",
X"FE0C",
X"02EE",
X"055F",
X"0A41",
X"0EA6",
X"0D2F",
X"09C4",
X"07D0",
X"03E8",
X"FE89",
X"FB9B",
X"F830",
X"F5BF",
X"F5BF",
X"FC18",
X"0000",
X"036B",
X"1117",
X"157C",
X"0F23",
X"FD8F",
X"FB1E",
X"FE0C",
X"F3CB",
X"EBFB",
X"F060",
X"F63C",
X"F2D1",
X"F92A",
X"01F4",
X"03E8",
X"07D0",
X"0D2F",
X"0E29",
X"0A41",
X"084D",
X"05DC",
X"0000",
X"FC95",
X"FAA1",
X"F736",
X"F542",
X"F8AD",
X"0000",
X"0177",
X"0BB8",
X"1676",
X"14FF",
X"05DC",
X"F830",
X"FD12",
X"F7B3",
X"EC78",
X"EB01",
X"F448",
X"F542",
X"F448",
X"FF06",
X"04E2",
X"0753",
X"0B3B",
X"0FA0",
X"0D2F",
X"09C4",
X"0659",
X"00FA",
X"FD12",
X"FB9B",
X"F92A",
X"F5BF",
X"F6B9",
X"FD8F",
X"01F4",
X"055F",
X"1405",
X"17ED",
X"0EA6",
X"FAA1",
X"F9A7",
X"FB1E",
X"EFE3",
X"E90D",
X"EF66",
X"F6B9",
X"F3CB",
X"FAA1",
X"0465",
X"05DC",
X"08CA",
X"0EA6",
X"0DAC",
X"084D",
X"05DC",
X"02EE",
X"FE0C",
X"FA24",
X"F92A",
X"F63C",
X"F736",
X"FB1E",
X"02EE",
X"02EE",
X"101D",
X"1A5E",
X"1405",
X"00FA",
X"F542",
X"FB1E",
X"F34E",
X"EA84",
X"EBFB",
X"F5BF",
X"F542",
X"F736",
X"0465",
X"084D",
X"07D0",
X"0D2F",
X"0F23",
X"09C4",
X"0659",
X"0465",
X"FF06",
X"FB1E",
X"FAA1",
X"F830",
X"F63C",
X"F8AD",
X"FF83",
X"03E8",
X"0B3B",
X"18E7",
X"157C",
X"0753",
X"F6B9",
X"F8AD",
X"F5BF",
X"EB01",
X"E98A",
X"F2D1",
X"F7B3",
X"F5BF",
X"007D",
X"0A41",
X"09C4",
X"0CB2",
X"0EA6",
X"0A41",
X"05DC",
X"04E2",
X"FF83",
X"FB1E",
X"FA24",
X"F8AD",
X"F736",
X"F9A7",
X"FE0C",
X"03E8",
X"08CA",
X"1676",
X"186A",
X"0CB2",
X"FAA1",
X"F34E",
X"F63C",
X"ED72",
X"E890",
X"ED72",
X"F736",
X"F8AD",
X"FC95",
X"08CA",
X"0ABE",
X"0B3B",
X"0F23",
X"0CB2",
X"06D6",
X"04E2",
X"00FA",
X"FB9B",
X"F9A7",
X"FA24",
X"F830",
X"F8AD",
X"FC95",
X"02EE",
X"07D0",
X"128E",
X"19E1",
X"101D",
X"0000",
X"F254",
X"F3CB",
X"EEE9",
X"E890",
X"EB7E",
X"F542",
X"FAA1",
X"FC18",
X"0659",
X"0C35",
X"0ABE",
X"0EA6",
X"0F23",
X"07D0",
X"02EE",
X"007D",
X"FC18",
X"FA24",
X"FB1E",
X"F92A",
X"F7B3",
X"FB9B",
X"00FA",
X"0659",
X"0DAC",
X"1964",
X"14FF",
X"055F",
X"F5BF",
X"F15A",
X"F060",
X"EA07",
X"E98A",
X"F15A",
X"FA24",
X"FD12",
X"0271",
X"0B3B",
X"0C35",
X"0C35",
X"0EA6",
X"0947",
X"036B",
X"0177",
X"FD8F",
X"F9A7",
X"FA24",
X"FB1E",
X"F92A",
X"FB1E",
X"0000",
X"055F",
X"0B3B",
X"16F3",
X"17ED",
X"0947",
X"F830",
X"EFE3",
X"EFE3",
X"EA07",
X"E890",
X"EEE9",
X"FA24",
X"FF83",
X"01F4",
X"09C4",
X"0D2F",
X"0D2F",
X"0EA6",
X"0A41",
X"036B",
X"FF83",
X"FE0C",
X"FAA1",
X"F9A7",
X"FB9B",
X"FAA1",
X"FB1E",
X"FF06",
X"02EE",
X"07D0",
X"1117",
X"1BD5",
X"1211",
X"0000",
X"F0DD",
X"ECF5",
X"EA84",
X"E796",
X"EB01",
X"F3CB",
X"FE89",
X"0271",
X"084D",
X"0FA0",
X"0E29",
X"0C35",
X"0CB2",
X"06D6",
X"FF83",
X"FD12",
X"FAA1",
X"F9A7",
X"FC18",
X"FC18",
X"FB1E",
X"FD8F",
X"01F4",
X"06D6",
X"0EA6",
X"1ADB",
X"16F3",
X"036B",
X"F1D7",
X"EA84",
X"EA84",
X"E796",
X"EA84",
X"F34E",
X"FF83",
X"05DC",
X"06D6",
X"0CB2",
X"0DAC",
X"0BB8",
X"0A41",
X"0465",
X"FE89",
X"FD12",
X"FC95",
X"FB1E",
X"FC18",
X"FE89",
X"FD12",
X"FD8F",
X"007D",
X"04E2",
X"08CA",
X"1482",
X"1C52",
X"0D2F",
X"F92A",
X"EA84",
X"E890",
X"E890",
X"EA84",
X"EF66",
X"FAA1",
X"055F",
X"0753",
X"0ABE",
X"0F23",
X"0BB8",
X"084D",
X"055F",
X"007D",
X"FC95",
X"FC18",
X"FAA1",
X"FB9B",
X"FE89",
X"FE89",
X"FD8F",
X"007D",
X"036B",
X"06D6",
X"0FA0",
X"1D4C",
X"1405",
X"FE89",
X"ECF5",
X"E69C",
X"E813",
X"E90D",
X"EE6C",
X"F736",
X"03E8",
X"0947",
X"0947",
X"0DAC",
X"0CB2",
X"0947",
X"055F",
X"FF83",
X"FB9B",
X"FD12",
X"FC18",
X"FB1E",
X"FD8F",
X"00FA",
X"0000",
X"FF83",
X"0177",
X"055F",
X"0CB2",
X"1964",
X"18E7",
X"04E2",
X"F15A",
X"E69C",
X"E5A2",
X"E813",
X"ED72",
X"F542",
X"01F4",
X"0BB8",
X"0BB8",
X"0CB2",
X"0E29",
X"084D",
X"03E8",
X"007D",
X"FB9B",
X"FA24",
X"FB1E",
X"FC18",
X"FE0C",
X"00FA",
X"00FA",
X"FF83",
X"0177",
X"03E8",
X"08CA",
X"128E",
X"1A5E",
X"0E29",
X"F92A",
X"EA84",
X"E525",
X"E719",
X"EB01",
X"F15A",
X"FB9B",
X"084D",
X"0C35",
X"0ABE",
X"0C35",
X"0ABE",
X"0659",
X"01F4",
X"FE0C",
X"FAA1",
X"FA24",
X"FC95",
X"FE0C",
X"00FA",
X"01F4",
X"0000",
X"007D",
X"0177",
X"055F",
X"0BB8",
X"19E1",
X"186A",
X"036B",
X"F15A",
X"E5A2",
X"E525",
X"E90D",
X"EFE3",
X"F63C",
X"01F4",
X"0CB2",
X"0BB8",
X"0ABE",
X"0BB8",
X"07D0",
X"02EE",
X"FE89",
X"FC18",
X"FAA1",
X"FB1E",
X"FC95",
X"FD8F",
X"0177",
X"0177",
X"0000",
X"01F4",
X"0465",
X"0A41",
X"157C",
X"1D4C",
X"0C35",
X"F6B9",
X"E890",
X"E3AE",
X"E719",
X"ED72",
X"F448",
X"FC18",
X"0947",
X"0EA6",
X"0ABE",
X"0ABE",
X"0947",
X"0465",
X"FE89",
X"FB1E",
X"FA24",
X"FC18",
X"FE89",
X"FF83",
X"01F4",
X"0271",
X"0000",
X"FF83",
X"007D",
X"055F",
X"0DAC",
X"1B58",
X"14FF",
X"FE89",
X"EDEF",
X"E331",
X"E4A8",
X"EBFB",
X"F448",
X"FA24",
X"04E2",
X"0EA6",
X"0C35",
X"0A41",
X"09C4",
X"055F",
X"0000",
X"FC18",
X"FB9B",
X"FC95",
X"FD8F",
X"FF83",
X"01F4",
X"036B",
X"007D",
X"FE0C",
X"FE89",
X"0177",
X"0753",
X"157C",
X"1DC9",
X"09C4",
X"F542",
X"E69C",
X"E2B4",
X"E98A",
X"F254",
X"F92A",
X"FE0C",
X"0A41",
X"0E29",
X"09C4",
X"09C4",
X"07D0",
X"0271",
X"FD12",
X"FB9B",
X"FC18",
X"FD12",
X"FE89",
X"FF83",
X"01F4",
X"0271",
X"0000",
X"FF83",
X"0177",
X"06D6",
X"128E",
X"1E46",
X"101D",
X"F830",
X"E90D",
X"E043",
X"E525",
X"EFE3",
X"F8AD",
X"FE0C",
X"084D",
X"0FA0",
X"0ABE",
X"06D6",
X"0659",
X"0465",
X"FF06",
X"FB9B",
X"FC95",
X"FE0C",
X"FF06",
X"FF83",
X"00FA",
X"0271",
X"0000",
X"FD8F",
X"FF06",
X"04E2",
X"0EA6",
X"1C52",
X"1770",
X"FF83",
X"EE6C",
X"E4A8",
X"E237",
X"EB01",
X"F5BF",
X"FD8F",
X"04E2",
X"0CB2",
X"0BB8",
X"06D6",
X"05DC",
X"04E2",
X"007D",
X"FC18",
X"FC18",
X"FD8F",
X"FF06",
X"007D",
X"0177",
X"0271",
X"0271",
X"FF06",
X"FF06",
X"036B",
X"09C4",
X"16F3",
X"19E1",
X"07D0",
X"F2D1",
X"E61F",
X"E0C0",
X"E719",
X"F3CB",
X"FAA1",
X"0177",
X"0A41",
X"0D2F",
X"0A41",
X"084D",
X"0753",
X"036B",
X"FE0C",
X"FB9B",
X"FD12",
X"FE89",
X"FF83",
X"0000",
X"0000",
X"00FA",
X"FF83",
X"FE0C",
X"00FA",
X"0659",
X"109A",
X"1B58",
X"128E",
X"FB9B",
X"EB7E",
X"E2B4",
X"E3AE",
X"EEE9",
X"F7B3",
X"FD8F",
X"055F",
X"0BB8",
X"0ABE",
X"0753",
X"06D6",
X"04E2",
X"00FA",
X"FC95",
X"FC95",
X"FF06",
X"FF06",
X"00FA",
X"01F4",
X"01F4",
X"00FA",
X"FE0C",
X"FD12",
X"007D",
X"08CA",
X"1676",
X"1C52",
X"09C4",
X"F2D1",
X"E719",
X"E13D",
X"E719",
X"F3CB",
X"FC18",
X"00FA",
X"08CA",
X"0DAC",
X"0A41",
X"07D0",
X"05DC",
X"02EE",
X"FE89",
X"FC18",
X"FE0C",
X"FF06",
X"007D",
X"0177",
X"01F4",
X"0271",
X"FF83",
X"FD12",
X"FF06",
X"0465",
X"0D2F",
X"1B58",
X"15F9",
X"FC95",
X"EBFB",
X"E331",
X"E1BA",
X"EDEF",
X"FB9B",
X"007D",
X"036B",
X"0BB8",
X"0BB8",
X"06D6",
X"055F",
X"02EE",
X"FF83",
X"FC18",
X"FD12",
X"0000",
X"01F4",
X"02EE",
X"036B",
X"02EE",
X"0000",
X"FD8F",
X"FC18",
X"0000",
X"07D0",
X"15F9",
X"203A",
X"0BB8",
X"F3CB",
X"E813",
X"E0C0",
X"E525",
X"F34E",
X"FE89",
X"007D",
X"0753",
X"0DAC",
X"09C4",
X"055F",
X"03E8",
X"036B",
X"FE89",
X"FB1E",
X"FE0C",
X"00FA",
X"01F4",
X"036B",
X"03E8",
X"007D",
X"FE0C",
X"FB9B",
X"FC18",
X"0465",
X"0DAC",
X"1FBD",
X"1B58",
X"FD12",
X"EB7E",
X"E0C0",
X"E0C0",
X"EBFB",
X"FB9B",
X"0177",
X"01F4",
X"0C35",
X"0CB2",
X"07D0",
X"03E8",
X"01F4",
X"00FA",
X"FB9B",
X"FB1E",
X"FF06",
X"01F4",
X"036B",
X"03E8",
X"0177",
X"007D",
X"FD8F",
X"FAA1",
X"0000",
X"06D6",
X"1405",
X"22AB",
X"0E29",
X"F3CB",
X"E719",
X"E0C0",
X"E5A2",
X"F34E",
X"0000",
X"0000",
X"055F",
X"0CB2",
X"09C4",
X"05DC",
X"0177",
X"00FA",
X"FE89",
X"FB9B",
X"FE0C",
X"0177",
X"0271",
X"0271",
X"0177",
X"FF06",
X"FC18",
X"FAA1",
X"FC18",
X"0465",
X"0D2F",
X"1EC3",
X"1FBD",
X"01F4",
X"ED72",
X"E237",
X"DF49",
X"E90D",
X"F9A7",
X"01F4",
X"0177",
X"0947",
X"0CB2",
X"084D",
X"055F",
X"01F4",
X"0177",
X"FE0C",
X"FAA1",
X"FE89",
X"0177",
X"0271",
X"03E8",
X"01F4",
X"FD8F",
X"FB1E",
X"F9A7",
X"FE89",
X"07D0",
X"130B",
X"2328",
X"1482",
X"F7B3",
X"E890",
X"DF49",
X"E2B4",
X"F1D7",
X"FF83",
X"0177",
X"03E8",
X"0BB8",
X"0A41",
X"0659",
X"0271",
X"007D",
X"0000",
X"FC18",
X"FD12",
X"007D",
X"0271",
X"02EE",
X"03E8",
X"007D",
X"FC18",
X"FAA1",
X"FB9B",
X"036B",
X"0CB2",
X"1ADB",
X"21B1",
X"08CA",
X"EFE3",
X"E2B4",
X"DDD2",
X"E69C",
X"F7B3",
X"01F4",
X"0271",
X"06D6",
X"0CB2",
X"0947",
X"055F",
X"00FA",
X"007D",
X"0000",
X"FC95",
X"FF06",
X"01F4",
X"02EE",
X"0271",
X"0177",
X"FE0C",
X"FB1E",
X"FA24",
X"FC95",
X"06D6",
X"0D2F",
X"1CCF",
X"1D4C",
X"007D",
X"EC78",
X"E3AE",
X"E237",
X"EBFB",
X"FC18",
X"02EE",
X"0000",
X"0659",
X"0ABE",
X"0753",
X"0465",
X"0000",
X"00FA",
X"FE89",
X"FD8F",
X"00FA",
X"036B",
X"0271",
X"00FA",
X"FF83",
X"FB9B",
X"FA24",
X"F9A7",
X"007D",
X"08CA",
X"109A",
X"2422",
X"1676",
X"F8AD",
X"E90D",
X"E043",
X"E2B4",
X"EFE3",
X"0000",
X"0000",
X"FF06",
X"0947",
X"0B3B",
X"084D",
X"036B",
X"00FA",
X"00FA",
X"FE0C",
X"FF06",
X"01F4",
X"02EE",
X"FF83",
X"FF06",
X"FE0C",
X"FD12",
X"FD12",
X"FF06",
X"06D6",
X"09C4",
X"16F3",
X"21B1",
X"084D",
X"EFE3",
X"E4A8",
X"E043",
X"E719",
X"F830",
X"03E8",
X"FF83",
X"00FA",
X"09C4",
X"0A41",
X"0753",
X"0271",
X"01F4",
X"0000",
X"FD12",
X"FE0C",
X"0271",
X"0271",
X"FF06",
X"FF83",
X"FD8F",
X"FC18",
X"FD8F",
X"00FA",
X"084D",
X"09C4",
X"1ADB",
X"1EC3",
X"007D",
X"EB7E",
X"E2B4",
X"E13D",
X"EB01",
X"FD12",
X"036B",
X"FD12",
X"03E8",
X"0CB2",
X"0B3B",
X"0659",
X"00FA",
X"00FA",
X"FE0C",
X"FC95",
X"FE0C",
X"0271",
X"01F4",
X"0000",
X"0000",
X"FD12",
X"FD12",
X"0000",
X"0465",
X"08CA",
X"0A41",
X"1BD5",
X"1770",
X"F9A7",
X"E90D",
X"E42B",
X"E719",
X"F0DD",
X"FF83",
X"00FA",
X"FB9B",
X"0659",
X"0DAC",
X"0947",
X"0271",
X"FD8F",
X"0177",
X"FF83",
X"FE89",
X"007D",
X"007D",
X"FE0C",
X"FE89",
X"FF83",
X"FE0C",
X"0000",
X"0271",
X"06D6",
X"0947",
X"0C35",
X"1B58",
X"0FA0",
X"F3CB",
X"E61F",
X"E2B4",
X"E890",
X"F6B9",
X"036B",
X"0000",
X"FE0C",
X"09C4",
X"0DAC",
X"0947",
X"0177",
X"FC95",
X"FF06",
X"FD8F",
X"FD8F",
X"0000",
X"FE0C",
X"FC18",
X"0000",
X"007D",
X"FF83",
X"03E8",
X"055F",
X"07D0",
X"07D0",
X"0E29",
X"186A",
X"0753",
X"F1D7",
X"E796",
X"E525",
X"EB01",
X"F92A",
X"01F4",
X"FE0C",
X"00FA",
X"0A41",
X"0BB8",
X"084D",
X"00FA",
X"FE0C",
X"FE89",
X"FD12",
X"FF83",
X"007D",
X"FE0C",
X"FC18",
X"FF06",
X"FF83",
X"0000",
X"036B",
X"0465",
X"06D6",
X"0753",
X"1194",
X"15F9",
X"0271",
X"F1D7",
X"E890",
X"E796",
X"EE6C",
X"FB1E",
X"00FA",
X"FE89",
X"0271",
X"0A41",
X"0ABE",
X"07D0",
X"01F4",
X"007D",
X"0000",
X"FF06",
X"007D",
X"FF83",
X"FC95",
X"FC18",
X"FF06",
X"FF83",
X"00FA",
X"03E8",
X"055F",
X"06D6",
X"07D0",
X"1211",
X"1211",
X"FF83",
X"F2D1",
X"EB01",
X"E98A",
X"F060",
X"FB9B",
X"FF83",
X"FE89",
X"0465",
X"0ABE",
X"0A41",
X"0659",
X"007D",
X"00FA",
X"FF06",
X"FE0C",
X"0000",
X"FF06",
X"FC95",
X"FD12",
X"FF06",
X"FE89",
X"00FA",
X"03E8",
X"05DC",
X"06D6",
X"06D6",
X"101D",
X"0D2F",
X"FD8F",
X"F4C5",
X"ED72",
X"EB7E",
X"F2D1",
X"FB9B",
X"FE89",
X"0000",
X"0659",
X"0A41",
X"084D",
X"03E8",
X"0000",
X"00FA",
X"FE89",
X"FE89",
X"FF06",
X"FE0C",
X"FC95",
X"FE0C",
X"FF06",
X"FF06",
X"01F4",
X"03E8",
X"055F",
X"05DC",
X"07D0",
X"0FA0",
X"0B3B",
X"FE89",
X"F5BF",
X"EFE3",
X"EF66",
X"F4C5",
X"FAA1",
X"FC95",
X"FE89",
X"05DC",
X"0A41",
X"0947",
X"03E8",
X"007D",
X"0000",
X"FE89",
X"FF06",
X"FE89",
X"FD8F",
X"FD8F",
X"007D",
X"00FA",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"02EE",
X"084D",
X"084D",
X"036B",
X"FF83",
X"FAA1",
X"F830",
X"F8AD",
X"F830",
X"F736",
X"F7B3",
X"FE89",
X"04E2",
X"0753",
X"06D6",
X"055F",
X"0465",
X"0271",
X"007D",
X"FE0C",
X"FB9B",
X"FB1E",
X"FE0C",
X"007D",
X"0177",
X"0271",
X"01F4",
X"007D",
X"0000",
X"007D",
X"0465",
X"03E8",
X"0271",
X"0177",
X"FE89",
X"FD12",
X"FB9B",
X"F92A",
X"F736",
X"F830",
X"FE0C",
X"02EE",
X"04E2",
X"055F",
X"055F",
X"04E2",
X"02EE",
X"0000",
X"FD8F",
X"FB1E",
X"FB9B",
X"FE89",
X"0000",
X"0177",
X"02EE",
X"02EE",
X"01F4",
X"00FA",
X"01F4",
X"03E8",
X"0271",
X"01F4",
X"0177",
X"FE89",
X"FD8F",
X"FB9B",
X"F9A7",
X"F7B3",
X"F9A7",
X"FF06",
X"0271",
X"03E8",
X"0465",
X"0465",
X"036B",
X"0177",
X"FF83",
X"FC95",
X"FB1E",
X"FD12",
X"FF83",
X"0177",
X"02EE",
X"036B",
X"02EE",
X"01F4",
X"00FA",
X"01F4",
X"0271",
X"00FA",
X"0177",
X"0000",
X"FE0C",
X"FD8F",
X"FB9B",
X"F9A7",
X"F8AD",
X"FB9B",
X"0000",
X"01F4",
X"036B",
X"03E8",
X"0465",
X"036B",
X"0177",
X"FF06",
X"FC18",
X"FB9B",
X"FD12",
X"FF83",
X"0177",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"02EE",
X"0177",
X"0000",
X"00FA",
X"FF83",
X"FE89",
X"FD8F",
X"FB1E",
X"F92A",
X"F92A",
X"FD12",
X"007D",
X"0271",
X"03E8",
X"03E8",
X"03E8",
X"02EE",
X"00FA",
X"FF06",
X"FC95",
X"FC95",
X"FE0C",
X"FF83",
X"0177",
X"0271",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"0000",
X"FF06",
X"FD12",
X"FB9B",
X"FC18",
X"FE89",
X"0000",
X"007D",
X"0177",
X"01F4",
X"01F4",
X"0177",
X"007D",
X"FF83",
X"FE0C",
X"FE89",
X"0000",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FF83",
X"FF06",
X"007D",
X"0177",
X"0177",
X"00FA",
X"FF06",
X"FD12",
X"FC18",
X"FD12",
X"FF06",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"0177",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FE89",
X"FF83",
X"0000",
X"0177",
X"0271",
X"0271",
X"01F4",
X"FF83",
X"FD12",
X"FC18",
X"FD12",
X"FE89",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"0177",
X"007D",
X"0000",
X"FF83",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FF83",
X"0000",
X"007D",
X"01F4",
X"01F4",
X"01F4",
X"00FA",
X"FF06",
X"FD12",
X"FC95",
X"FD8F",
X"FF06",
X"FF06",
X"FF06",
X"0000",
X"007D",
X"00FA",
X"0177",
X"00FA",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF06",
X"FF06",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"01F4",
X"0177",
X"007D",
X"FE89",
X"FD12",
X"FD12",
X"FE89",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"00FA",
X"0177",
X"0177",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"FF83",
X"FE0C",
X"FD8F",
X"FE89",
X"0000",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"00FA",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"FF06",
X"FE89",
X"FE89",
X"FF83",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"007D",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"0177",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FF06",
X"FF83",
X"007D",
X"007D",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FD8F",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"007D",
X"0177",
X"0177",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD12",
X"FC95",
X"FC18",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"00FA",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0177",
X"007D",
X"FF83",
X"FE0C",
X"FD12",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FD8F",
X"FE89",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"0000",
X"0000",
X"00FA",
X"0177",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"0177",
X"0000",
X"FE89",
X"FD12",
X"FC18",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FE0C",
X"FF06",
X"007D",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"00FA",
X"FF83",
X"FE0C",
X"FC95",
X"FB9B",
X"FB1E",
X"FB1E",
X"FB9B",
X"FD12",
X"FE0C",
X"FF83",
X"00FA",
X"01F4",
X"02EE",
X"02EE",
X"02EE",
X"01F4",
X"0177",
X"007D",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"0177",
X"0271",
X"02EE",
X"036B",
X"036B",
X"0271",
X"00FA",
X"FF06",
X"FD12",
X"FB9B",
X"FAA1",
X"FAA1",
X"FAA1",
X"FB9B",
X"FD12",
X"FF06",
X"007D",
X"01F4",
X"02EE",
X"036B",
X"036B",
X"02EE",
X"01F4",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"007D",
X"01F4",
X"02EE",
X"036B",
X"036B",
X"036B",
X"01F4",
X"007D",
X"FE89",
X"FC95",
X"FB1E",
X"FAA1",
X"FAA1",
X"FB1E",
X"FC18",
X"FD8F",
X"FF06",
X"007D",
X"01F4",
X"02EE",
X"036B",
X"02EE",
X"0271",
X"0177",
X"007D",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"0271",
X"036B",
X"03E8",
X"03E8",
X"02EE",
X"01F4",
X"0000",
X"FE0C",
X"FC18",
X"FB1E",
X"FA24",
X"FA24",
X"FB1E",
X"FC95",
X"FE0C",
X"FF83",
X"00FA",
X"0271",
X"02EE",
X"036B",
X"02EE",
X"0271",
X"0177",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"02EE",
X"03E8",
X"03E8",
X"03E8",
X"02EE",
X"0177",
X"FF83",
X"FD12",
X"FB9B",
X"FA24",
X"F9A7",
X"FA24",
X"FB1E",
X"FD12",
X"FE89",
X"007D",
X"01F4",
X"02EE",
X"036B",
X"036B",
X"02EE",
X"01F4",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"00FA",
X"01F4",
X"036B",
X"03E8",
X"0465",
X"036B",
X"0271",
X"00FA",
X"FF06",
X"FC95",
X"FB1E",
X"F9A7",
X"F9A7",
X"F9A7",
X"FB1E",
X"FD12",
X"FF06",
X"007D",
X"0271",
X"036B",
X"03E8",
X"036B",
X"02EE",
X"01F4",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FF06",
X"FF83",
X"00FA",
X"01F4",
X"036B",
X"0465",
X"0465",
X"03E8",
X"0271",
X"00FA",
X"FE89",
X"FC95",
X"FAA1",
X"F9A7",
X"F92A",
X"F9A7",
X"FB1E",
X"FD12",
X"FF06",
X"00FA",
X"0271",
X"036B",
X"03E8",
X"03E8",
X"036B",
X"0271",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FF83",
X"007D",
X"01F4",
X"036B",
X"0465",
X"0465",
X"03E8",
X"0271",
X"00FA",
X"FE89",
X"FC18",
X"FA24",
X"F92A",
X"F92A",
X"F9A7",
X"FB1E",
X"FD12",
X"FF06",
X"00FA",
X"0271",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"01F4",
X"00FA",
X"FF83",
X"FE89",
X"FE89",
X"FE89",
X"FF83",
X"00FA",
X"0271",
X"03E8",
X"04E2",
X"04E2",
X"03E8",
X"0271",
X"007D",
X"FE89",
X"FB9B",
X"F9A7",
X"F92A",
X"F8AD",
X"F9A7",
X"FB1E",
X"FD8F",
X"FF83",
X"0177",
X"02EE",
X"03E8",
X"0465",
X"03E8",
X"02EE",
X"01F4",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FE89",
X"FF83",
X"00FA",
X"02EE",
X"03E8",
X"04E2",
X"04E2",
X"03E8",
X"0271",
X"007D",
X"FE0C",
X"FB1E",
X"F9A7",
X"F8AD",
X"F8AD",
X"F9A7",
X"FB9B",
X"FD8F",
X"0000",
X"0177",
X"036B",
X"03E8",
X"0465",
X"03E8",
X"02EE",
X"01F4",
X"007D",
X"FF83",
X"FE89",
X"FE89",
X"FF06",
X"0000",
X"0177",
X"02EE",
X"0465",
X"055F",
X"04E2",
X"03E8",
X"01F4",
X"0000",
X"FD8F",
X"FAA1",
X"F92A",
X"F830",
X"F830",
X"F92A",
X"FB9B",
X"FD8F",
X"0000",
X"01F4",
X"036B",
X"0465",
X"0465",
X"03E8",
X"02EE",
X"01F4",
X"007D",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"0000",
X"01F4",
X"036B",
X"04E2",
X"055F",
X"04E2",
X"03E8",
X"01F4",
X"0000",
X"FD12",
X"FAA1",
X"F8AD",
X"F830",
X"F830",
X"F92A",
X"FB9B",
X"FD8F",
X"0000",
X"01F4",
X"036B",
X"0465",
X"0465",
X"03E8",
X"02EE",
X"01F4",
X"007D",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"0000",
X"01F4",
X"036B",
X"04E2",
X"055F",
X"04E2",
X"036B",
X"01F4",
X"FF83",
X"FD12",
X"FA24",
X"F8AD",
X"F830",
X"F830",
X"F9A7",
X"FB9B",
X"FE0C",
X"0000",
X"01F4",
X"036B",
X"0465",
X"0465",
X"03E8",
X"02EE",
X"01F4",
X"007D",
X"FF06",
X"FE0C",
X"FE0C",
X"FE89",
X"0000",
X"01F4",
X"03E8",
X"04E2",
X"055F",
X"04E2",
X"036B",
X"0177",
X"FF83",
X"FC95",
X"FA24",
X"F8AD",
X"F7B3",
X"F830",
X"F9A7",
X"FC18",
X"FE89",
X"007D",
X"0271",
X"03E8",
X"0465",
X"0465",
X"03E8",
X"02EE",
X"0177",
X"0000",
X"FF06",
X"FE0C",
X"FE89",
X"FF06",
X"007D",
X"0271",
X"03E8",
X"055F",
X"05DC",
X"04E2",
X"036B",
X"0177",
X"FF06",
X"FC18",
X"F9A7",
X"F830",
X"F7B3",
X"F830",
X"F9A7",
X"FC18",
X"FE89",
X"007D",
X"0271",
X"03E8",
X"0465",
X"0465",
X"03E8",
X"02EE",
X"0177",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FF83",
X"007D",
X"0271",
X"03E8",
X"04E2",
X"055F",
X"04E2",
X"036B",
X"0177",
X"FF06",
X"FC18",
X"F9A7",
X"F830",
X"F7B3",
X"F830",
X"F9A7",
X"FC18",
X"FE89",
X"007D",
X"0271",
X"03E8",
X"0465",
X"0465",
X"03E8",
X"02EE",
X"0177",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"007D",
X"01F4",
X"03E8",
X"04E2",
X"055F",
X"0465",
X"036B",
X"0177",
X"FF06",
X"FC18",
X"F9A7",
X"F830",
X"F7B3",
X"F830",
X"F9A7",
X"FC18",
X"FE89",
X"007D",
X"0271",
X"03E8",
X"04E2",
X"04E2",
X"0465",
X"02EE",
X"01F4",
X"007D",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"007D",
X"0271",
X"03E8",
X"04E2",
X"055F",
X"0465",
X"036B",
X"0177",
X"FF06",
X"FB9B",
X"F92A",
X"F830",
X"F7B3",
X"F830",
X"F9A7",
X"FC18",
X"FE89",
X"007D",
X"0271",
X"0465",
X"04E2",
X"04E2",
X"0465",
X"036B",
X"01F4",
X"007D",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"007D",
X"01F4",
X"03E8",
X"04E2",
X"055F",
X"0465",
X"036B",
X"0177",
X"FE89",
X"FB9B",
X"F92A",
X"F830",
X"F7B3",
X"F830",
X"F9A7",
X"FC18",
X"FE89",
X"007D",
X"0271",
X"0465",
X"04E2",
X"04E2",
X"0465",
X"036B",
X"01F4",
X"007D",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"007D",
X"01F4",
X"03E8",
X"04E2",
X"04E2",
X"0465",
X"036B",
X"0177",
X"FE89",
X"FB9B",
X"F9A7",
X"F830",
X"F7B3",
X"F830",
X"F9A7",
X"FC18",
X"FE0C",
X"007D",
X"02EE",
X"0465",
X"04E2",
X"04E2",
X"04E2",
X"036B",
X"01F4",
X"007D",
X"FF06",
X"FE89",
X"FE0C",
X"FF06",
X"007D",
X"01F4",
X"03E8",
X"04E2",
X"055F",
X"04E2",
X"036B",
X"0177",
X"FE89",
X"FB9B",
X"F92A",
X"F7B3",
X"F736",
X"F7B3",
X"F9A7",
X"FC18",
X"FE89",
X"00FA",
X"02EE",
X"0465",
X"055F",
X"055F",
X"04E2",
X"036B",
X"01F4",
X"0000",
X"FE89",
X"FE0C",
X"FE0C",
X"FF06",
X"007D",
X"0271",
X"0465",
X"055F",
X"055F",
X"04E2",
X"036B",
X"00FA",
X"FE0C",
X"FB1E",
X"F8AD",
X"F7B3",
X"F736",
X"F7B3",
X"F9A7",
X"FC18",
X"FE89",
X"00FA",
X"036B",
X"04E2",
X"055F",
X"055F",
X"04E2",
X"036B",
X"01F4",
X"0000",
X"FE89",
X"FE0C",
X"FE0C",
X"FF06",
X"007D",
X"0271",
X"0465",
X"055F",
X"055F",
X"04E2",
X"036B",
X"00FA",
X"FE0C",
X"FB1E",
X"F92A",
X"F7B3",
X"F736",
X"F7B3",
X"F9A7",
X"FC18",
X"FE89",
X"00FA",
X"036B",
X"04E2",
X"055F",
X"055F",
X"04E2",
X"036B",
X"01F4",
X"0000",
X"FE89",
X"FE0C",
X"FD8F",
X"FE89",
X"0000",
X"01F4",
X"03E8",
X"055F",
X"05DC",
X"055F",
X"03E8",
X"00FA",
X"FE0C",
X"FB1E",
X"F92A",
X"F7B3",
X"F6B9",
X"F7B3",
X"F92A",
X"FB9B",
X"FE89",
X"00FA",
X"036B",
X"04E2",
X"05DC",
X"05DC",
X"055F",
X"03E8",
X"01F4",
X"0000",
X"FE89",
X"FD8F",
X"FD8F",
X"FE89",
X"0000",
X"0271",
X"0465",
X"055F",
X"05DC",
X"055F",
X"036B",
X"00FA",
X"FE0C",
X"FAA1",
X"F8AD",
X"F736",
X"F6B9",
X"F736",
X"F92A",
X"FB9B",
X"FE89",
X"00FA",
X"036B",
X"055F",
X"0659",
X"0659",
X"055F",
X"03E8",
X"01F4",
X"0000",
X"FE89",
X"FD8F",
X"FD8F",
X"FE89",
X"007D",
X"0271",
X"04E2",
X"0659",
X"0659",
X"055F",
X"03E8",
X"00FA",
X"FD8F",
X"FAA1",
X"F830",
X"F6B9",
X"F63C",
X"F6B9",
X"F8AD",
X"FB1E",
X"FE0C",
X"00FA",
X"03E8",
X"055F",
X"0659",
X"0659",
X"05DC",
X"03E8",
X"01F4",
X"0000",
X"FE0C",
X"FD12",
X"FD8F",
X"FE89",
X"0000",
X"0271",
X"04E2",
X"0659",
X"06D6",
X"0659",
X"03E8",
X"00FA",
X"FD8F",
X"FAA1",
X"F830",
X"F63C",
X"F5BF",
X"F6B9",
X"F8AD",
X"FB1E",
X"FE0C",
X"0177",
X"03E8",
X"055F",
X"0659",
X"0659",
X"055F",
X"03E8",
X"01F4",
X"0000",
X"FE0C",
X"FD12",
X"FD12",
X"FE0C",
X"0000",
X"0271",
X"04E2",
X"06D6",
X"0753",
X"0659",
X"0465",
X"0177",
X"FE0C",
X"FAA1",
X"F830",
X"F5BF",
X"F542",
X"F5BF",
X"F830",
X"FAA1",
X"FE0C",
X"00FA",
X"03E8",
X"05DC",
X"0753",
X"0753",
X"0659",
X"04E2",
X"0271",
X"0000",
X"FE0C",
X"FC95",
X"FC95",
X"FE0C",
X"FF83",
X"0271",
X"04E2",
X"06D6",
X"07D0",
X"06D6",
X"0465",
X"0177",
X"FE0C",
X"FAA1",
X"F7B3",
X"F542",
X"F4C5",
X"F542",
X"F7B3",
X"FAA1",
X"FE0C",
X"0177",
X"0465",
X"0659",
X"07D0",
X"07D0",
X"06D6",
X"04E2",
X"02EE",
X"0000",
X"FD8F",
X"FC18",
X"FC18",
X"FD12",
X"FF06",
X"01F4",
X"0465",
X"06D6",
X"07D0",
X"0753",
X"055F",
X"01F4",
X"FE89",
X"FAA1",
X"F736",
X"F4C5",
X"F3CB",
X"F4C5",
X"F736",
X"FA24",
X"FD8F",
X"00FA",
X"0465",
X"06D6",
X"07D0",
X"07D0",
X"06D6",
X"055F",
X"02EE",
X"0000",
X"FD8F",
X"FC18",
X"FB9B",
X"FC95",
X"FE89",
X"0177",
X"0465",
X"0753",
X"0947",
X"08CA",
X"06D6",
X"036B",
X"FF83",
X"FB1E",
X"F736",
X"F3CB",
X"F2D1",
X"F3CB",
X"F63C",
X"F9A7",
X"FD8F",
X"0177",
X"04E2",
X"07D0",
X"0947",
X"08CA",
X"07D0",
X"05DC",
X"02EE",
X"0000",
X"FD12",
X"FB9B",
X"FB1E",
X"FC18",
X"FE0C",
X"00FA",
X"0465",
X"0753",
X"0947",
X"0947",
X"06D6",
X"036B",
X"FF83",
X"FAA1",
X"F6B9",
X"F34E",
X"F254",
X"F2D1",
X"F5BF",
X"F92A",
X"FD12",
X"0177",
X"04E2",
X"07D0",
X"0947",
X"0947",
X"084D",
X"0659",
X"03E8",
X"007D",
X"FD8F",
X"FB9B",
X"FAA1",
X"FB1E",
X"FD12",
X"0000",
X"036B",
X"0753",
X"09C4",
X"0A41",
X"084D",
X"04E2",
X"007D",
X"FB1E",
X"F63C",
X"F254",
X"F0DD",
X"F15A",
X"F448",
X"F7B3",
X"FC95",
X"00FA",
X"055F",
X"084D",
X"0A41",
X"0A41",
X"0947",
X"06D6",
X"03E8",
X"007D",
X"FD12",
X"FAA1",
X"F9A7",
X"FA24",
X"FC95",
X"0000",
X"03E8",
X"07D0",
X"0ABE",
X"0BB8",
X"09C4",
X"0659",
X"0177",
X"FB9B",
X"F63C",
X"F1D7",
X"F060",
X"F0DD",
X"F3CB",
X"F7B3",
X"FC18",
X"00FA",
X"04E2",
X"084D",
X"0A41",
X"0A41",
X"0947",
X"0753",
X"03E8",
X"007D",
X"FD12",
X"FAA1",
X"F9A7",
X"FA24",
X"FC18",
X"FF83",
X"036B",
X"07D0",
X"0B3B",
X"0CB2",
X"0B3B",
X"07D0",
X"0271",
X"FC18",
X"F5BF",
X"F15A",
X"EF66",
X"EFE3",
X"F254",
X"F6B9",
X"FB9B",
X"00FA",
X"055F",
X"08CA",
X"0ABE",
X"0ABE",
X"09C4",
X"0753",
X"0465",
X"00FA",
X"FD8F",
X"FB1E",
X"F9A7",
X"FA24",
X"FB9B",
X"FE89",
X"0271",
X"06D6",
X"0ABE",
X"0CB2",
X"0C35",
X"08CA",
X"02EE",
X"FC18",
X"F5BF",
X"F15A",
X"EEE9",
X"EF66",
X"F1D7",
X"F5BF",
X"FAA1",
X"0000",
X"0465",
X"084D",
X"0A41",
X"0ABE",
X"09C4",
X"07D0",
X"0465",
X"00FA",
X"FE0C",
X"FB1E",
X"F92A",
X"F9A7",
X"FB1E",
X"FE0C",
X"0177",
X"0659",
X"0ABE",
X"0D2F",
X"0CB2",
X"0947",
X"036B",
X"FC95",
X"F5BF",
X"F0DD",
X"EE6C",
X"EE6C",
X"F15A",
X"F5BF",
X"FB1E",
X"007D",
X"05DC",
X"09C4",
X"0BB8",
X"0BB8",
X"0ABE",
X"084D",
X"0465",
X"00FA",
X"FD12",
X"FA24",
X"F8AD",
X"F92A",
X"FAA1",
X"FD8F",
X"00FA",
X"055F",
X"09C4",
X"0D2F",
X"0DAC",
X"0ABE",
X"03E8",
X"FC95",
X"F542",
X"F060",
X"EDEF",
X"EDEF",
X"F0DD",
X"F5BF",
X"FB9B",
X"00FA",
X"05DC",
X"09C4",
X"0B3B",
X"0B3B",
X"0A41",
X"07D0",
X"0465",
X"007D",
X"FD12",
X"FAA1",
X"F8AD",
X"F8AD",
X"FA24",
X"FD12",
X"00FA",
X"05DC",
X"0ABE",
X"0E29",
X"0F23",
X"0BB8",
X"0465",
X"FB9B",
X"F448",
X"EEE9",
X"EC78",
X"ECF5",
X"F060",
X"F5BF",
X"FB9B",
X"0177",
X"0659",
X"09C4",
X"0BB8",
X"0C35",
X"0ABE",
X"07D0",
X"0465",
X"00FA",
X"FE0C",
X"FB1E",
X"F92A",
X"F92A",
X"FAA1",
X"FD8F",
X"01F4",
X"0659",
X"0ABE",
X"0F23",
X"101D",
X"0C35",
X"036B",
X"FAA1",
X"F34E",
X"EE6C",
X"EB7E",
X"EC78",
X"F060",
X"F5BF",
X"FC18",
X"0271",
X"0753",
X"0ABE",
X"0C35",
X"0C35",
X"0ABE",
X"0753",
X"036B",
X"0000",
X"FC95",
X"FA24",
X"F8AD",
X"F8AD",
X"FAA1",
X"FE0C",
X"0271",
X"06D6",
X"0BB8",
X"101D",
X"109A",
X"0BB8",
X"01F4",
X"F8AD",
X"F1D7",
X"ECF5",
X"EA84",
X"EC78",
X"F0DD",
X"F6B9",
X"FD8F",
X"0465",
X"0947",
X"0BB8",
X"0D2F",
X"0CB2",
X"09C4",
X"05DC",
X"01F4",
X"FE0C",
X"FB9B",
X"F9A7",
X"F92A",
X"F9A7",
X"FC18",
X"0000",
X"03E8",
X"084D",
X"0D2F",
X"1194",
X"1211",
X"0BB8",
X"00FA",
X"F6B9",
X"F060",
X"EB7E",
X"E90D",
X"EB01",
X"F060",
X"F736",
X"FE89",
X"05DC",
X"0A41",
X"0CB2",
X"0E29",
X"0CB2",
X"0947",
X"04E2",
X"007D",
X"FD12",
X"FAA1",
X"F9A7",
X"F92A",
X"FAA1",
X"FD8F",
X"01F4",
X"055F",
X"08CA",
X"0DAC",
X"1211",
X"1194",
X"0947",
X"FD12",
X"F34E",
X"EE6C",
X"EA07",
X"E90D",
X"EBFB",
X"F2D1",
X"FA24",
X"0177",
X"084D",
X"0BB8",
X"0DAC",
X"0DAC",
X"0BB8",
X"0753",
X"0271",
X"FE0C",
X"FB9B",
X"FA24",
X"FA24",
X"FAA1",
X"FC18",
X"FF83",
X"036B",
X"0659",
X"09C4",
X"0E29",
X"1211",
X"1117",
X"0753",
X"FA24",
X"F1D7",
X"ECF5",
X"E90D",
X"E890",
X"ED72",
X"F4C5",
X"FC18",
X"03E8",
X"09C4",
X"0C35",
X"0D2F",
X"0CB2",
X"0A41",
X"05DC",
X"00FA",
X"FD12",
X"FB1E",
X"F9A7",
X"F92A",
X"F9A7",
X"FC18",
X"0000",
X"03E8",
X"07D0",
X"0BB8",
X"1117",
X"1388",
X"0F23",
X"036B",
X"F6B9",
X"EFE3",
X"EBFB",
X"E98A",
X"EA84",
X"F0DD",
X"F8AD",
X"FF83",
X"06D6",
X"0B3B",
X"0C35",
X"0CB2",
X"0B3B",
X"07D0",
X"02EE",
X"FF06",
X"FB9B",
X"FA24",
X"F9A7",
X"F9A7",
X"FB1E",
X"FE0C",
X"01F4",
X"05DC",
X"0A41",
X"0E29",
X"130B",
X"130B",
X"0B3B",
X"FC95",
X"F0DD",
X"EB7E",
X"E890",
X"E796",
X"EB7E",
X"F448",
X"FC95",
X"03E8",
X"0A41",
X"0D2F",
X"0D2F",
X"0D2F",
X"0ABE",
X"0659",
X"0177",
X"FC95",
X"FA24",
X"F9A7",
X"F9A7",
X"FA24",
X"FC95",
X"007D",
X"055F",
X"08CA",
X"0CB2",
X"101D",
X"130B",
X"0FA0",
X"055F",
X"F63C",
X"EBFB",
X"E90D",
X"E796",
X"E813",
X"ED72",
X"F736",
X"007D",
X"07D0",
X"0D2F",
X"0E29",
X"0DAC",
X"0C35",
X"084D",
X"02EE",
X"FD8F",
X"FAA1",
X"F92A",
X"FA24",
X"FAA1",
X"FC95",
X"FF83",
X"036B",
X"07D0",
X"0B3B",
X"0EA6",
X"1211",
X"130B",
X"0CB2",
X"FF06",
X"F060",
X"E90D",
X"E719",
X"E61F",
X"E90D",
X"F15A",
X"FC18",
X"03E8",
X"0B3B",
X"0F23",
X"0EA6",
X"0D2F",
X"0ABE",
X"05DC",
X"007D",
X"FC18",
X"F9A7",
X"F9A7",
X"FA24",
X"FB9B",
X"FE0C",
X"0177",
X"04E2",
X"08CA",
X"0C35",
X"0F23",
X"130B",
X"1211",
X"08CA",
X"F9A7",
X"EBFB",
X"E796",
X"E69C",
X"E61F",
X"EA84",
X"F5BF",
X"00FA",
X"07D0",
X"0DAC",
X"0FA0",
X"0DAC",
X"0BB8",
X"0753",
X"0271",
X"FD8F",
X"FA24",
X"F92A",
X"FAA1",
X"FC18",
X"FD8F",
X"0000",
X"0271",
X"05DC",
X"0947",
X"0CB2",
X"109A",
X"1405",
X"109A",
X"04E2",
X"F4C5",
X"E890",
X"E525",
X"E525",
X"E69C",
X"ED72",
X"F9A7",
X"0465",
X"0C35",
X"109A",
X"101D",
X"0DAC",
X"0A41",
X"04E2",
X"FF06",
X"FAA1",
X"F830",
X"F8AD",
X"FAA1",
X"FC18",
X"FE0C",
X"00FA",
X"0465",
X"0753",
X"0ABE",
X"0EA6",
X"130B",
X"157C",
X"0EA6",
X"FF83",
X"EE6C",
X"E525",
X"E42B",
X"E42B",
X"E813",
X"F254",
X"0000",
X"0947",
X"0EA6",
X"1194",
X"0F23",
X"0B3B",
X"06D6",
X"0177",
X"FC18",
X"F8AD",
X"F830",
X"FA24",
X"FC95",
X"FE0C",
X"0000",
X"02EE",
X"05DC",
X"08CA",
X"0BB8",
X"0FA0",
X"1482",
X"1482",
X"09C4",
X"F8AD",
X"EA07",
X"E42B",
X"E42B",
X"E5A2",
X"EB7E",
X"F7B3",
X"0465",
X"0BB8",
X"101D",
X"109A",
X"0CB2",
X"08CA",
X"0465",
X"FE0C",
X"F9A7",
X"F830",
X"F8AD",
X"FB9B",
X"FD8F",
X"FF06",
X"0177",
X"0465",
X"06D6",
X"08CA",
X"0C35",
X"1117",
X"1676",
X"1388",
X"0465",
X"F254",
X"E69C",
X"E3AE",
X"E3AE",
X"E719",
X"EFE3",
X"FD12",
X"07D0",
X"0DAC",
X"109A",
X"0FA0",
X"0ABE",
X"0659",
X"0177",
X"FC95",
X"F92A",
X"F8AD",
X"FA24",
X"FC95",
X"FE89",
X"007D",
X"036B",
X"055F",
X"06D6",
X"09C4",
X"0EA6",
X"1388",
X"16F3",
X"0E29",
X"FB9B",
X"EA84",
X"E331",
X"E331",
X"E5A2",
X"EA07",
X"F4C5",
X"0271",
X"0C35",
X"101D",
X"1117",
X"0DAC",
X"08CA",
X"0465",
X"FF06",
X"FA24",
X"F7B3",
X"F7B3",
X"F9A7",
X"FD12",
X"FF06",
X"0177",
X"03E8",
X"0659",
X"08CA",
X"0B3B",
X"0F23",
X"1405",
X"157C",
X"09C4",
X"F7B3",
X"E890",
X"E3AE",
X"E42B",
X"E69C",
X"EBFB",
X"F830",
X"0659",
X"0E29",
X"109A",
X"109A",
X"0D2F",
X"08CA",
X"02EE",
X"FD8F",
X"F92A",
X"F7B3",
X"F92A",
X"FC18",
X"FE0C",
X"FF06",
X"00FA",
X"036B",
X"0659",
X"0947",
X"0DAC",
X"1405",
X"1964",
X"130B",
X"0000",
X"ED72",
X"E3AE",
X"E237",
X"E3AE",
X"E719",
X"F0DD",
X"FF83",
X"0A41",
X"0EA6",
X"101D",
X"0F23",
X"0A41",
X"055F",
X"0000",
X"FB1E",
X"F8AD",
X"F92A",
X"FB9B",
X"FE0C",
X"FF06",
X"0000",
X"01F4",
X"03E8",
X"05DC",
X"07D0",
X"0BB8",
X"1388",
X"1964",
X"1117",
X"FC95",
X"EA07",
X"E13D",
X"E13D",
X"E4A8",
X"E98A",
X"F4C5",
X"036B",
X"0D2F",
X"109A",
X"109A",
X"0DAC",
X"084D",
X"036B",
X"FE0C",
X"F92A",
X"F830",
X"FA24",
X"FC95",
X"FF06",
X"0000",
X"00FA",
X"0271",
X"0465",
X"0659",
X"0947",
X"0E29",
X"15F9",
X"1ADB",
X"0F23",
X"F92A",
X"E719",
X"DFC6",
X"E13D",
X"E525",
X"EC78",
X"F830",
X"07D0",
X"109A",
X"1194",
X"0FA0",
X"0BB8",
X"04E2",
X"FF06",
X"FB9B",
X"F9A7",
X"F9A7",
X"FB9B",
X"FF06",
X"00FA",
X"01F4",
X"00FA",
X"007D",
X"02EE",
X"055F",
X"084D",
X"0E29",
X"186A",
X"1C52",
X"0BB8",
X"F34E",
X"E1BA",
X"DC5B",
X"E043",
X"E719",
X"EF66",
X"FD12",
X"0C35",
X"1211",
X"0FA0",
X"0D2F",
X"08CA",
X"02EE",
X"FE89",
X"FAA1",
X"F92A",
X"FA24",
X"FD8F",
X"0177",
X"0271",
X"0271",
X"01F4",
X"0271",
X"03E8",
X"04E2",
X"084D",
X"0E29",
X"186A",
X"1BD5",
X"08CA",
X"F060",
X"E13D",
X"DECC",
X"E3AE",
X"EB01",
X"F2D1",
X"FF06",
X"0D2F",
X"109A",
X"0DAC",
X"0ABE",
X"0659",
X"00FA",
X"FD12",
X"FA24",
X"FA24",
X"FB9B",
X"FF06",
X"02EE",
X"03E8",
X"036B",
X"0271",
X"01F4",
X"0271",
X"03E8",
X"08CA",
X"101D",
X"1CCF",
X"1BD5",
X"036B",
X"EB7E",
X"DDD2",
X"DDD2",
X"E525",
X"EE6C",
X"F6B9",
X"02EE",
X"0FA0",
X"1117",
X"0D2F",
X"0947",
X"02EE",
X"FD12",
X"FB1E",
X"FAA1",
X"FAA1",
X"FC95",
X"00FA",
X"036B",
X"036B",
X"02EE",
X"01F4",
X"00FA",
X"007D",
X"036B",
X"08CA",
X"0FA0",
X"1BD5",
X"1BD5",
X"036B",
X"EB7E",
X"DD55",
X"DE4F",
X"E61F",
X"EE6C",
X"F5BF",
X"0271",
X"1194",
X"130B",
X"0D2F",
X"084D",
X"036B",
X"FD8F",
X"FA24",
X"F9A7",
X"FAA1",
X"FD12",
X"0271",
X"05DC",
X"04E2",
X"02EE",
X"007D",
X"FF83",
X"007D",
X"03E8",
X"0B3B",
X"130B",
X"1F40",
X"18E7",
X"FD12",
X"E61F",
X"DC5B",
X"DFC6",
X"E813",
X"F254",
X"FAA1",
X"0659",
X"128E",
X"1194",
X"0ABE",
X"0659",
X"0177",
X"FC18",
X"F92A",
X"F92A",
X"FAA1",
X"FE89",
X"02EE",
X"06D6",
X"05DC",
X"03E8",
X"00FA",
X"FE89",
X"007D",
X"036B",
X"08CA",
X"0F23",
X"1D4C",
X"1BD5",
X"FF83",
X"E796",
X"DC5B",
X"DF49",
X"E719",
X"F1D7",
X"FB1E",
X"05DC",
X"1211",
X"109A",
X"084D",
X"02EE",
X"FF06",
X"FB1E",
X"F9A7",
X"FB1E",
X"FD12",
X"00FA",
X"055F",
X"0753",
X"0465",
X"01F4",
X"0000",
X"FD12",
X"FE89",
X"00FA",
X"05DC",
X"0DAC",
X"1E46",
X"2134",
X"02EE",
X"E813",
X"DBDE",
X"DE4F",
X"E69C",
X"F1D7",
X"FC95",
X"03E8",
X"109A",
X"1117",
X"09C4",
X"0465",
X"FF83",
X"FB1E",
X"F830",
X"FB1E",
X"FE89",
X"0271",
X"055F",
X"05DC",
X"02EE",
X"0177",
X"0000",
X"FC95",
X"FE0C",
X"007D",
X"05DC",
X"0E29",
X"1EC3",
X"23A5",
X"055F",
X"E90D",
X"DBDE",
X"DDD2",
X"E5A2",
X"F15A",
X"FC18",
X"0271",
X"1117",
X"130B",
X"0A41",
X"0177",
X"FC18",
X"F92A",
X"F7B3",
X"FB9B",
X"0000",
X"04E2",
X"0753",
X"06D6",
X"0465",
X"0177",
X"FF06",
X"FB9B",
X"FF83",
X"01F4",
X"0659",
X"0C35",
X"1BD5",
X"23A5",
X"055F",
X"E890",
X"DBDE",
X"DE4F",
X"E813",
X"F542",
X"00FA",
X"036B",
X"0E29",
X"0FA0",
X"0753",
X"0000",
X"FA24",
X"F830",
X"F7B3",
X"FC95",
X"01F4",
X"0659",
X"0753",
X"084D",
X"0659",
X"02EE",
X"0000",
X"FB1E",
X"FC95",
X"0000",
X"03E8",
X"0753",
X"17ED",
X"2616",
X"09C4",
X"EA07",
X"DBDE",
X"DE4F",
X"E98A",
X"F6B9",
X"01F4",
X"02EE",
X"0BB8",
X"0FA0",
X"0659",
X"FD8F",
X"F92A",
X"FA24",
X"F9A7",
X"FD12",
X"01F4",
X"06D6",
X"0947",
X"09C4",
X"06D6",
X"01F4",
X"FF06",
X"FB1E",
X"FB1E",
X"FD12",
X"0177",
X"0753",
X"17ED",
X"280A",
X"0EA6",
X"EC78",
X"DD55",
X"DDD2",
X"E719",
X"F448",
X"0177",
X"036B",
X"0A41",
X"0F23",
X"0753",
X"FF83",
X"FAA1",
X"FAA1",
X"F92A",
X"FB1E",
X"00FA",
X"06D6",
X"08CA",
X"08CA",
X"06D6",
X"00FA",
X"FE89",
X"FB1E",
X"FAA1",
X"FC95",
X"00FA",
X"0659",
X"130B",
X"2693",
X"157C",
X"F2D1",
X"E1BA",
X"DECC",
X"E61F",
X"F254",
X"FF83",
X"0271",
X"0753",
X"0F23",
X"0947",
X"0177",
X"FB9B",
X"FC18",
X"FB1E",
X"FB1E",
X"FF83",
X"0465",
X"08CA",
X"084D",
X"0659",
X"0000",
X"FE0C",
X"FC95",
X"F9A7",
X"FAA1",
X"007D",
X"0659",
X"109A",
X"249F",
X"19E1",
X"F63C",
X"E237",
X"DECC",
X"E4A8",
X"F060",
X"0000",
X"055F",
X"06D6",
X"0EA6",
X"0B3B",
X"0177",
X"FB9B",
X"FB1E",
X"FAA1",
X"F9A7",
X"FF83",
X"036B",
X"084D",
X"0947",
X"06D6",
X"007D",
X"FE89",
X"FD8F",
X"F9A7",
X"FB1E",
X"0000",
X"04E2",
X"0ABE",
X"203A",
X"1FBD",
X"FD8F",
X"E61F",
X"E043",
X"E42B",
X"ECF5",
X"FC18",
X"0465",
X"036B",
X"0B3B",
X"0C35",
X"036B",
X"FD12",
X"FC18",
X"FE89",
X"FC95",
X"FF83",
X"01F4",
X"06D6",
X"0947",
X"0753",
X"007D",
X"FD12",
X"FC95",
X"F830",
X"F92A",
X"FE89",
X"05DC",
X"0ABE",
X"1D4C",
X"249F",
X"04E2",
X"E813",
X"E0C0",
X"E331",
X"E98A",
X"F830",
X"04E2",
X"036B",
X"084D",
X"0DAC",
X"05DC",
X"FD8F",
X"FAA1",
X"FE0C",
X"FC95",
X"0000",
X"02EE",
X"0659",
X"0947",
X"0753",
X"01F4",
X"FD12",
X"FD12",
X"F830",
X"F736",
X"FC18",
X"02EE",
X"084D",
X"17ED",
X"2887",
X"0FA0",
X"EDEF",
X"E13D",
X"E237",
X"E69C",
X"F2D1",
X"0271",
X"02EE",
X"05DC",
X"0EA6",
X"08CA",
X"FE0C",
X"F92A",
X"FE0C",
X"FE89",
X"0000",
X"02EE",
X"055F",
X"0947",
X"07D0",
X"0271",
X"FC18",
X"FD8F",
X"F9A7",
X"F63C",
X"FAA1",
X"01F4",
X"07D0",
X"1388",
X"280A",
X"17ED",
X"F34E",
X"E2B4",
X"E237",
X"E5A2",
X"F060",
X"0177",
X"0465",
X"036B",
X"0ABE",
X"084D",
X"FF83",
X"F9A7",
X"FD12",
X"0000",
X"0177",
X"0465",
X"055F",
X"084D",
X"07D0",
X"036B",
X"FC95",
X"FC95",
X"FC18",
X"F736",
X"FA24",
X"00FA",
X"06D6",
X"0E29",
X"222E",
X"1EC3",
X"FB9B",
X"E5A2",
X"E331",
X"E61F",
X"EDEF",
X"FD12",
X"036B",
X"00FA",
X"0753",
X"084D",
X"0177",
X"FB9B",
X"FD12",
X"0177",
X"01F4",
X"036B",
X"036B",
X"06D6",
X"07D0",
X"055F",
X"FD8F",
X"FAA1",
X"FC95",
X"F9A7",
X"F9A7",
X"FF06",
X"05DC",
X"0A41",
X"1ADB",
X"2422",
X"0659",
X"EB7E",
X"E42B",
X"E525",
X"EA84",
X"F7B3",
X"01F4",
X"FF83",
X"04E2",
X"09C4",
X"0465",
X"FE89",
X"FD12",
X"00FA",
X"00FA",
X"02EE",
X"02EE",
X"0465",
X"0753",
X"0753",
X"00FA",
X"FA24",
X"FC95",
X"FB1E",
X"F9A7",
X"FD12",
X"02EE",
X"0753",
X"1482",
X"2693",
X"128E",
X"F15A",
X"E3AE",
X"E331",
X"E890",
X"F448",
X"00FA",
X"0177",
X"036B",
X"09C4",
X"05DC",
X"FF83",
X"FC95",
X"FF06",
X"0000",
X"01F4",
X"0271",
X"036B",
X"0753",
X"084D",
X"036B",
X"FB1E",
X"FB9B",
X"FC18",
X"FA24",
X"FC18",
X"0177",
X"06D6",
X"0EA6",
X"2328",
X"1B58",
X"F8AD",
X"E525",
X"E237",
X"E61F",
X"F060",
X"FF83",
X"036B",
X"0271",
X"0947",
X"08CA",
X"01F4",
X"FD12",
X"FD8F",
X"FF06",
X"0000",
X"0271",
X"0177",
X"04E2",
X"07D0",
X"04E2",
X"FC95",
X"FB1E",
X"FE0C",
X"FC18",
X"FC95",
X"007D",
X"05DC",
X"09C4",
X"1C52",
X"21B1",
X"01F4",
X"E813",
X"E331",
X"E61F",
X"ED72",
X"FC18",
X"02EE",
X"007D",
X"05DC",
X"09C4",
X"036B",
X"FE0C",
X"FE0C",
X"FF83",
X"007D",
X"02EE",
X"01F4",
X"03E8",
X"06D6",
X"0659",
X"FE0C",
X"FA24",
X"FE0C",
X"FD12",
X"FC18",
X"FD8F",
X"0271",
X"06D6",
X"1482",
X"251C",
X"0F23",
X"EEE9",
X"E4A8",
X"E69C",
X"EB01",
X"F5BF",
X"00FA",
X"FF83",
X"01F4",
X"09C4",
X"0659",
X"007D",
X"FF06",
X"007D",
X"FF83",
X"0000",
X"00FA",
X"02EE",
X"084D",
X"0947",
X"0177",
X"F9A7",
X"FC95",
X"FD12",
X"FB1E",
X"FB9B",
X"FF83",
X"0465",
X"0CB2",
X"222E",
X"1ADB",
X"F92A",
X"E796",
X"E61F",
X"E98A",
X"F0DD",
X"FE0C",
X"0177",
X"FF83",
X"0753",
X"084D",
X"01F4",
X"FF06",
X"00FA",
X"00FA",
X"FF83",
X"00FA",
X"01F4",
X"06D6",
X"09C4",
X"03E8",
X"FB1E",
X"FB1E",
X"FD12",
X"FAA1",
X"FAA1",
X"FD8F",
X"03E8",
X"09C4",
X"1B58",
X"222E",
X"04E2",
X"EB01",
X"E525",
X"E890",
X"EDEF",
X"FA24",
X"02EE",
X"FF06",
X"036B",
X"08CA",
X"0465",
X"FF83",
X"FF83",
X"007D",
X"FF06",
X"0000",
X"01F4",
X"05DC",
X"0A41",
X"06D6",
X"FE0C",
X"FA24",
X"FB9B",
X"FAA1",
X"FA24",
X"FC95",
X"01F4",
X"0753",
X"130B",
X"23A5",
X"1211",
X"F254",
X"E61F",
X"E796",
X"EC78",
X"F542",
X"0000",
X"FF83",
X"0000",
X"0753",
X"06D6",
X"0177",
X"FF83",
X"00FA",
X"007D",
X"FF83",
X"0177",
X"03E8",
X"08CA",
X"07D0",
X"00FA",
X"FB1E",
X"FB9B",
X"FB9B",
X"F9A7",
X"FAA1",
X"FF83",
X"05DC",
X"0D2F",
X"1F40",
X"1C52",
X"FC95",
X"E90D",
X"E719",
X"EB01",
X"F15A",
X"FC18",
X"FF83",
X"FE89",
X"0465",
X"0753",
X"03E8",
X"007D",
X"007D",
X"01F4",
X"007D",
X"0000",
X"0177",
X"0659",
X"0947",
X"04E2",
X"FE0C",
X"FB1E",
X"FB1E",
X"F8AD",
X"F92A",
X"FD12",
X"036B",
X"09C4",
X"18E7",
X"21B1",
X"0947",
X"EDEF",
X"E61F",
X"E90D",
X"EF66",
X"F92A",
X"FF83",
X"FE89",
X"01F4",
X"0753",
X"05DC",
X"00FA",
X"FE89",
X"007D",
X"0177",
X"00FA",
X"00FA",
X"03E8",
X"08CA",
X"0659",
X"0000",
X"FB9B",
X"FB9B",
X"FA24",
X"F92A",
X"FC18",
X"007D",
X"0659",
X"1211",
X"222E",
X"157C",
X"F830",
X"E796",
X"E525",
X"EB01",
X"F448",
X"FD8F",
X"FF83",
X"00FA",
X"07D0",
X"07D0",
X"02EE",
X"FF06",
X"FF83",
X"0177",
X"0177",
X"007D",
X"007D",
X"05DC",
X"0753",
X"02EE",
X"FE89",
X"FD12",
X"FB1E",
X"F8AD",
X"FAA1",
X"FE0C",
X"03E8",
X"0CB2",
X"1E46",
X"1CCF",
X"00FA",
X"EB7E",
X"E4A8",
X"E98A",
X"F15A",
X"FA24",
X"FE0C",
X"FE89",
X"055F",
X"0947",
X"0659",
X"0177",
X"FF83",
X"00FA",
X"0177",
X"0177",
X"FF83",
X"03E8",
X"0753",
X"0465",
X"FF83",
X"FD12",
X"FB9B",
X"F92A",
X"FAA1",
X"FC95",
X"0271",
X"09C4",
X"18E7",
X"1F40",
X"08CA",
X"EF66",
X"E4A8",
X"E796",
X"EF66",
X"F92A",
X"FF06",
X"FE89",
X"03E8",
X"08CA",
X"06D6",
X"0271",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"007D",
X"036B",
X"0753",
X"05DC",
X"007D",
X"FC95",
X"FB1E",
X"F8AD",
X"F9A7",
X"FC18",
X"01F4",
X"084D",
X"1482",
X"1F40",
X"0F23",
X"F4C5",
X"E61F",
X"E61F",
X"ECF5",
X"F63C",
X"FF06",
X"FF06",
X"0271",
X"084D",
X"07D0",
X"0465",
X"007D",
X"FF83",
X"FF83",
X"00FA",
X"00FA",
X"01F4",
X"055F",
X"0659",
X"0271",
X"FE0C",
X"FC95",
X"F92A",
X"F9A7",
X"FC18",
X"0177",
X"0753",
X"0F23",
X"1C52",
X"1388",
X"FB9B",
X"EA84",
X"E5A2",
X"EB01",
X"F3CB",
X"FE89",
X"FF83",
X"00FA",
X"0753",
X"06D6",
X"03E8",
X"0177",
X"FF83",
X"FE89",
X"0000",
X"0177",
X"0177",
X"04E2",
X"06D6",
X"03E8",
X"FF83",
X"FD12",
X"FA24",
X"F9A7",
X"FC95",
X"00FA",
X"0659",
X"0CB2",
X"17ED",
X"14FF",
X"0000",
X"EF66",
X"E719",
X"E98A",
X"F1D7",
X"FC18",
X"007D",
X"0177",
X"06D6",
X"06D6",
X"03E8",
X"0177",
X"0000",
X"FF06",
X"FF83",
X"0177",
X"01F4",
X"0465",
X"05DC",
X"03E8",
X"0000",
X"FD12",
X"FB1E",
X"F9A7",
X"FC95",
X"00FA",
X"0659",
X"0B3B",
X"1405",
X"1405",
X"02EE",
X"F34E",
X"E98A",
X"E890",
X"EEE9",
X"F92A",
X"0000",
X"01F4",
X"06D6",
X"07D0",
X"0465",
X"0271",
X"007D",
X"FF83",
X"FF06",
X"007D",
X"007D",
X"02EE",
X"05DC",
X"04E2",
X"01F4",
X"FF83",
X"FE89",
X"FC95",
X"FD8F",
X"0000",
X"0465",
X"07D0",
X"0DAC",
X"101D",
X"0465",
X"F7B3",
X"EE6C",
X"EB01",
X"EF66",
X"F7B3",
X"FF06",
X"007D",
X"0465",
X"05DC",
X"036B",
X"0271",
X"01F4",
X"00FA",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"03E8",
X"03E8",
X"01F4",
X"FF83",
X"FF06",
X"FE0C",
X"FE89",
X"00FA",
X"0465",
X"0753",
X"09C4",
X"0C35",
X"04E2",
X"FB1E",
X"F34E",
X"EE6C",
X"EFE3",
X"F5BF",
X"FD8F",
X"00FA",
X"0465",
X"055F",
X"0271",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0177",
X"0271",
X"036B",
X"036B",
X"00FA",
X"0000",
X"FF83",
X"FF83",
X"00FA",
X"0271",
X"03E8",
X"055F",
X"084D",
X"03E8",
X"FC18",
X"F63C",
X"F1D7",
X"F254",
X"F5BF",
X"FB1E",
X"FE89",
X"01F4",
X"0465",
X"036B",
X"0271",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"02EE",
X"0465",
X"0465",
X"0177",
X"FF83",
X"FE0C",
X"FC18",
X"FB9B",
X"FC95",
X"FF06",
X"00FA",
X"036B",
X"0659",
X"04E2",
X"036B",
X"0177",
X"FE89",
X"FD12",
X"FB1E",
X"F8AD",
X"F63C",
X"F7B3",
X"FB1E",
X"FE89",
X"0271",
X"04E2",
X"0659",
X"06D6",
X"0659",
X"0465",
X"01F4",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FD12",
X"FE0C",
X"FF83",
X"01F4",
X"04E2",
X"055F",
X"04E2",
X"036B",
X"007D",
X"FE0C",
X"FB9B",
X"F8AD",
X"F63C",
X"F7B3",
X"F9A7",
X"FD12",
X"0177",
X"0465",
X"0659",
X"06D6",
X"05DC",
X"03E8",
X"01F4",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"0000",
X"0271",
X"036B",
X"03E8",
X"036B",
X"0177",
X"FF83",
X"FD12",
X"FAA1",
X"F7B3",
X"F736",
X"F8AD",
X"FB1E",
X"FF06",
X"0271",
X"04E2",
X"05DC",
X"05DC",
X"04E2",
X"036B",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"FF83",
X"FE89",
X"FE0C",
X"FD8F",
X"FE0C",
X"FF06",
X"00FA",
X"0271",
X"036B",
X"02EE",
X"0177",
X"FF06",
X"FC95",
X"FAA1",
X"F92A",
X"F8AD",
X"F9A7",
X"FB9B",
X"FF83",
X"0271",
X"0465",
X"055F",
X"04E2",
X"0465",
X"036B",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FE89",
X"FD12",
X"FD12",
X"FD8F",
X"FF83",
X"007D",
X"0177",
X"0271",
X"02EE",
X"0271",
X"0000",
X"FC95",
X"FA24",
X"F92A",
X"F92A",
X"FAA1",
X"FC95",
X"0000",
X"02EE",
X"04E2",
X"055F",
X"04E2",
X"0465",
X"036B",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"FF83",
X"FE0C",
X"FC95",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"01F4",
X"036B",
X"036B",
X"0271",
X"0000",
X"FE0C",
X"FD12",
X"FC18",
X"FB9B",
X"FB9B",
X"FD12",
X"FF83",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"00FA",
X"FE89",
X"FC18",
X"FB9B",
X"FC18",
X"FD12",
X"FE0C",
X"FE89",
X"00FA",
X"02EE",
X"03E8",
X"036B",
X"00FA",
X"FF06",
X"FE0C",
X"FC95",
X"FC18",
X"FB9B",
X"FD12",
X"FF06",
X"007D",
X"0177",
X"0271",
X"02EE",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0177",
X"FF83",
X"FD12",
X"FC18",
X"FC18",
X"FD12",
X"FE0C",
X"FE89",
X"0000",
X"0271",
X"03E8",
X"036B",
X"01F4",
X"FF83",
X"FE89",
X"FD12",
X"FC18",
X"FB9B",
X"FC18",
X"FE0C",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"036B",
X"036B",
X"0271",
X"01F4",
X"0000",
X"FD8F",
X"FC18",
X"FC18",
X"FC95",
X"FE0C",
X"FE89",
X"0000",
X"01F4",
X"036B",
X"036B",
X"0271",
X"0000",
X"FE89",
X"FD8F",
X"FC95",
X"FB9B",
X"FC18",
X"FD8F",
X"FF83",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"007D",
X"FE89",
X"FD12",
X"FC95",
X"FD8F",
X"FE89",
X"FE89",
X"FF06",
X"007D",
X"01F4",
X"0271",
X"01F4",
X"007D",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FC95",
X"FD8F",
X"FF06",
X"0000",
X"007D",
X"0177",
X"01F4",
X"02EE",
X"036B",
X"036B",
X"036B",
X"02EE",
X"01F4",
X"00FA",
X"FF06",
X"FD12",
X"FC95",
X"FC95",
X"FD8F",
X"FD8F",
X"FE0C",
X"FF83",
X"00FA",
X"01F4",
X"01F4",
X"00FA",
X"0000",
X"0000",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FF83",
X"0000",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0271",
X"01F4",
X"0177",
X"0000",
X"FE89",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"0271",
X"01F4",
X"0177",
X"007D",
X"FF06",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"0000",
X"007D",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0000",
X"FF06",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FF83",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF06",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"007D",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"007D",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"0271",
X"0271",
X"0271",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FC95",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"0271",
X"0271",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FD8F",
X"FD12",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"0177",
X"01F4",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FC18",
X"FC95",
X"FD8F",
X"FE89",
X"0000",
X"00FA",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"007D",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"00FA",
X"0000",
X"FF06",
X"FD8F",
X"FC95",
X"FC18",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FE0C",
X"FF06",
X"007D",
X"0177",
X"0271",
X"02EE",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"007D",
X"0177",
X"01F4",
X"0271",
X"0271",
X"01F4",
X"0177",
X"0000",
X"FE89",
X"FD8F",
X"FC18",
X"FB9B",
X"FB1E",
X"FB1E",
X"FB9B",
X"FC95",
X"FE0C",
X"FF83",
X"007D",
X"01F4",
X"02EE",
X"036B",
X"036B",
X"02EE",
X"0271",
X"0177",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"0271",
X"0271",
X"02EE",
X"0271",
X"0177",
X"0000",
X"FE89",
X"FD12",
X"FB9B",
X"FAA1",
X"FAA1",
X"FAA1",
X"FB9B",
X"FD12",
X"FE89",
X"0000",
X"0177",
X"02EE",
X"036B",
X"03E8",
X"03E8",
X"036B",
X"0271",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"01F4",
X"0271",
X"02EE",
X"0271",
X"01F4",
X"00FA",
X"FF83",
X"FE0C",
X"FC95",
X"FB9B",
X"FAA1",
X"FAA1",
X"FB1E",
X"FC18",
X"FD12",
X"FF06",
X"007D",
X"01F4",
X"02EE",
X"03E8",
X"03E8",
X"03E8",
X"02EE",
X"01F4",
X"007D",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"01F4",
X"0271",
X"02EE",
X"0271",
X"01F4",
X"00FA",
X"FF83",
X"FD8F",
X"FC18",
X"FB1E",
X"FAA1",
X"FAA1",
X"FB1E",
X"FC18",
X"FD8F",
X"FF06",
X"00FA",
X"0271",
X"036B",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0177",
X"007D",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"007D",
X"FF06",
X"FD8F",
X"FC18",
X"FAA1",
X"FA24",
X"FAA1",
X"FB1E",
X"FC95",
X"FE0C",
X"FF83",
X"0177",
X"02EE",
X"03E8",
X"0465",
X"03E8",
X"036B",
X"0271",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"0177",
X"007D",
X"FE89",
X"FD12",
X"FB9B",
X"FAA1",
X"FA24",
X"FAA1",
X"FB9B",
X"FC95",
X"FE89",
X"0000",
X"01F4",
X"036B",
X"0465",
X"0465",
X"03E8",
X"036B",
X"01F4",
X"007D",
X"FF83",
X"FE89",
X"FE89",
X"FE89",
X"FF83",
X"007D",
X"01F4",
X"02EE",
X"036B",
X"036B",
X"02EE",
X"01F4",
X"0000",
X"FE0C",
X"FC95",
X"FB1E",
X"FA24",
X"F9A7",
X"FAA1",
X"FB9B",
X"FD12",
X"FE89",
X"007D",
X"0271",
X"03E8",
X"0465",
X"04E2",
X"03E8",
X"02EE",
X"01F4",
X"007D",
X"FF06",
X"FE89",
X"FE0C",
X"FE89",
X"FF83",
X"00FA",
X"0271",
X"036B",
X"036B",
X"036B",
X"0271",
X"0177",
X"0000",
X"FE0C",
X"FC18",
X"FB1E",
X"FA24",
X"F9A7",
X"FA24",
X"FB9B",
X"FD12",
X"FF06",
X"00FA",
X"02EE",
X"0465",
X"04E2",
X"04E2",
X"03E8",
X"02EE",
X"0177",
X"0000",
X"FE89",
X"FE0C",
X"FD8F",
X"FE89",
X"FF83",
X"00FA",
X"0271",
X"036B",
X"03E8",
X"036B",
X"02EE",
X"01F4",
X"0000",
X"FE0C",
X"FC18",
X"FAA1",
X"F9A7",
X"F9A7",
X"FA24",
X"FB9B",
X"FD12",
X"FF06",
X"0177",
X"036B",
X"0465",
X"055F",
X"04E2",
X"0465",
X"02EE",
X"00FA",
X"FF83",
X"FE0C",
X"FD8F",
X"FD12",
X"FE0C",
X"FF83",
X"00FA",
X"02EE",
X"03E8",
X"0465",
X"03E8",
X"036B",
X"01F4",
X"0000",
X"FE0C",
X"FB9B",
X"FA24",
X"F9A7",
X"F92A",
X"FA24",
X"FB9B",
X"FD12",
X"FF83",
X"0177",
X"036B",
X"0465",
X"055F",
X"04E2",
X"03E8",
X"0271",
X"00FA",
X"FF06",
X"FE0C",
X"FD12",
X"FD12",
X"FE0C",
X"FF83",
X"0177",
X"036B",
X"0465",
X"04E2",
X"0465",
X"036B",
X"0271",
X"007D",
X"FE0C",
X"FB9B",
X"FA24",
X"F92A",
X"F92A",
X"F9A7",
X"FB1E",
X"FD12",
X"FF06",
X"0177",
X"036B",
X"04E2",
X"055F",
X"055F",
X"0465",
X"0271",
X"00FA",
X"FF06",
X"FD8F",
X"FD12",
X"FD12",
X"FE0C",
X"FF83",
X"0177",
X"036B",
X"0465",
X"04E2",
X"0465",
X"03E8",
X"0271",
X"007D",
X"FE0C",
X"FB9B",
X"FA24",
X"F92A",
X"F8AD",
X"F92A",
X"FB1E",
X"FC95",
X"FF06",
X"0177",
X"036B",
X"04E2",
X"055F",
X"055F",
X"0465",
X"0271",
X"007D",
X"FF06",
X"FD8F",
X"FC95",
X"FC95",
X"FD8F",
X"FF83",
X"0177",
X"036B",
X"04E2",
X"055F",
X"04E2",
X"0465",
X"02EE",
X"00FA",
X"FE0C",
X"FC18",
X"FA24",
X"F8AD",
X"F8AD",
X"F92A",
X"FAA1",
X"FC95",
X"FF06",
X"0177",
X"036B",
X"04E2",
X"05DC",
X"055F",
X"0465",
X"02EE",
X"00FA",
X"FF06",
X"FD12",
X"FC95",
X"FC95",
X"FD8F",
X"FF06",
X"00FA",
X"036B",
X"04E2",
X"055F",
X"055F",
X"04E2",
X"036B",
X"00FA",
X"FE89",
X"FC18",
X"FA24",
X"F8AD",
X"F830",
X"F8AD",
X"FA24",
X"FC18",
X"FE89",
X"0177",
X"036B",
X"04E2",
X"05DC",
X"05DC",
X"0465",
X"02EE",
X"00FA",
X"FF06",
X"FD12",
X"FC18",
X"FC95",
X"FD12",
X"FF06",
X"00FA",
X"036B",
X"04E2",
X"055F",
X"055F",
X"04E2",
X"036B",
X"00FA",
X"FE89",
X"FC18",
X"FA24",
X"F8AD",
X"F830",
X"F8AD",
X"FA24",
X"FC18",
X"FE89",
X"00FA",
X"036B",
X"04E2",
X"05DC",
X"05DC",
X"04E2",
X"02EE",
X"00FA",
X"FF06",
X"FD12",
X"FC18",
X"FC18",
X"FD12",
X"FE89",
X"00FA",
X"036B",
X"04E2",
X"05DC",
X"05DC",
X"04E2",
X"036B",
X"0177",
X"FF06",
X"FC95",
X"FAA1",
X"F92A",
X"F830",
X"F8AD",
X"F9A7",
X"FB9B",
X"FE0C",
X"00FA",
X"02EE",
X"04E2",
X"05DC",
X"05DC",
X"04E2",
X"036B",
X"00FA",
X"FF06",
X"FD12",
X"FC18",
X"FC18",
X"FC95",
X"FE89",
X"007D",
X"036B",
X"04E2",
X"05DC",
X"05DC",
X"055F",
X"0465",
X"01F4",
X"FF83",
X"FC95",
X"FAA1",
X"F8AD",
X"F7B3",
X"F7B3",
X"F92A",
X"FB1E",
X"FD8F",
X"007D",
X"02EE",
X"04E2",
X"05DC",
X"0659",
X"055F",
X"03E8",
X"01F4",
X"FF83",
X"FD8F",
X"FC18",
X"FB9B",
X"FC18",
X"FD8F",
X"0000",
X"0271",
X"04E2",
X"05DC",
X"0659",
X"0659",
X"04E2",
X"02EE",
X"007D",
X"FD8F",
X"FB1E",
X"F92A",
X"F7B3",
X"F736",
X"F830",
X"FA24",
X"FC95",
X"FF83",
X"0271",
X"04E2",
X"05DC",
X"0659",
X"05DC",
X"0465",
X"01F4",
X"0000",
X"FD8F",
X"FC18",
X"FB1E",
X"FB9B",
X"FD12",
X"FF83",
X"01F4",
X"04E2",
X"0659",
X"06D6",
X"06D6",
X"05DC",
X"036B",
X"00FA",
X"FE0C",
X"FB1E",
X"F92A",
X"F736",
X"F6B9",
X"F7B3",
X"F9A7",
X"FC18",
X"FF06",
X"01F4",
X"0465",
X"0659",
X"06D6",
X"0659",
X"04E2",
X"02EE",
X"007D",
X"FE0C",
X"FC18",
X"FB1E",
X"FB1E",
X"FC95",
X"FF06",
X"0177",
X"0465",
X"0659",
X"0753",
X"06D6",
X"05DC",
X"03E8",
X"00FA",
X"FE0C",
X"FB9B",
X"F92A",
X"F736",
X"F63C",
X"F736",
X"F92A",
X"FB9B",
X"FF06",
X"01F4",
X"04E2",
X"0659",
X"0753",
X"06D6",
X"055F",
X"02EE",
X"007D",
X"FD8F",
X"FB9B",
X"FAA1",
X"FAA1",
X"FC18",
X"FE89",
X"0177",
X"0465",
X"0659",
X"07D0",
X"0753",
X"0659",
X"0465",
X"01F4",
X"FF06",
X"FC18",
X"F92A",
X"F736",
X"F63C",
X"F6B9",
X"F8AD",
X"FB1E",
X"FE89",
X"0177",
X"0465",
X"0659",
X"0753",
X"0753",
X"05DC",
X"036B",
X"00FA",
X"FE0C",
X"FC18",
X"FAA1",
X"FAA1",
X"FB9B",
X"FD8F",
X"007D",
X"03E8",
X"0659",
X"07D0",
X"07D0",
X"06D6",
X"04E2",
X"0271",
X"FF83",
X"FC95",
X"F9A7",
X"F736",
X"F63C",
X"F63C",
X"F830",
X"FAA1",
X"FD8F",
X"00FA",
X"03E8",
X"0659",
X"0753",
X"0753",
X"05DC",
X"03E8",
X"0177",
X"FE89",
X"FC18",
X"FAA1",
X"FA24",
X"FB1E",
X"FD8F",
X"0000",
X"036B",
X"05DC",
X"07D0",
X"07D0",
X"0753",
X"055F",
X"02EE",
X"0000",
X"FD12",
X"FAA1",
X"F830",
X"F63C",
X"F63C",
X"F7B3",
X"F9A7",
X"FC95",
X"0000",
X"02EE",
X"055F",
X"06D6",
X"0753",
X"0659",
X"04E2",
X"0271",
X"FF83",
X"FD12",
X"FB1E",
X"FAA1",
X"FB1E",
X"FC95",
X"FF06",
X"01F4",
X"04E2",
X"06D6",
X"07D0",
X"07D0",
X"0659",
X"03E8",
X"00FA",
X"FE0C",
X"FB1E",
X"F8AD",
X"F6B9",
X"F63C",
X"F736",
X"F92A",
X"FB9B",
X"FF06",
X"01F4",
X"0465",
X"0659",
X"06D6",
X"0659",
X"04E2",
X"02EE",
X"007D",
X"FE0C",
X"FC18",
X"FB1E",
X"FB1E",
X"FC95",
X"FE89",
X"0177",
X"0465",
X"06D6",
X"07D0",
X"0753",
X"0659",
X"03E8",
X"0177",
X"FE89",
X"FC18",
X"F92A",
X"F736",
X"F63C",
X"F736",
X"F8AD",
X"FB1E",
X"FE0C",
X"00FA",
X"03E8",
X"05DC",
X"06D6",
X"0659",
X"055F",
X"036B",
X"00FA",
X"FE89",
X"FC95",
X"FB9B",
X"FB9B",
X"FC95",
X"FE89",
X"00FA",
X"03E8",
X"05DC",
X"06D6",
X"06D6",
X"05DC",
X"0465",
X"01F4",
X"FF83",
X"FC95",
X"FA24",
X"F830",
X"F6B9",
X"F6B9",
X"F830",
X"FA24",
X"FD12",
X"0000",
X"02EE",
X"055F",
X"0659",
X"06D6",
X"05DC",
X"03E8",
X"01F4",
X"FF83",
X"FD12",
X"FB9B",
X"FB1E",
X"FC18",
X"FE0C",
X"007D",
X"036B",
X"05DC",
X"0753",
X"0753",
X"0659",
X"04E2",
X"0271",
X"0000",
X"FD8F",
X"FAA1",
X"F830",
X"F63C",
X"F63C",
X"F7B3",
X"F9A7",
X"FC95",
X"FF83",
X"0271",
X"04E2",
X"0659",
X"06D6",
X"0659",
X"04E2",
X"0271",
X"0000",
X"FD8F",
X"FB9B",
X"FB1E",
X"FB9B",
X"FD12",
X"FF83",
X"0271",
X"04E2",
X"06D6",
X"07D0",
X"0753",
X"05DC",
X"036B",
X"00FA",
X"FE0C",
X"FB1E",
X"F830",
X"F63C",
X"F5BF",
X"F6B9",
X"F92A",
X"FB9B",
X"FF06",
X"01F4",
X"04E2",
X"06D6",
X"0753",
X"06D6",
X"055F",
X"02EE",
X"007D",
X"FE0C",
X"FC18",
X"FB1E",
X"FB1E",
X"FC95",
X"FE89",
X"01F4",
X"04E2",
X"06D6",
X"07D0",
X"07D0",
X"0659",
X"03E8",
X"0177",
X"FE89",
X"FB9B",
X"F8AD",
X"F63C",
X"F5BF",
X"F63C",
X"F830",
X"FB1E",
X"FE89",
X"01F4",
X"04E2",
X"06D6",
X"0753",
X"0753",
X"05DC",
X"036B",
X"00FA",
X"FE89",
X"FC18",
X"FAA1",
X"FAA1",
X"FB9B",
X"FD8F",
X"007D",
X"03E8",
X"06D6",
X"084D",
X"08CA",
X"07D0",
X"055F",
X"0271",
X"FF06",
X"FB9B",
X"F830",
X"F5BF",
X"F448",
X"F542",
X"F736",
X"FA24",
X"FE0C",
X"01F4",
X"04E2",
X"0753",
X"084D",
X"084D",
X"06D6",
X"0465",
X"0177",
X"FE89",
X"FB9B",
X"FA24",
X"F9A7",
X"FA24",
X"FC95",
X"FF83",
X"036B",
X"0659",
X"08CA",
X"0947",
X"08CA",
X"06D6",
X"036B",
X"0000",
X"FC18",
X"F8AD",
X"F5BF",
X"F3CB",
X"F448",
X"F63C",
X"F92A",
X"FD12",
X"00FA",
X"04E2",
X"0753",
X"08CA",
X"08CA",
X"07D0",
X"055F",
X"0271",
X"FF06",
X"FC18",
X"FA24",
X"F92A",
X"F92A",
X"FB1E",
X"FE89",
X"0271",
X"05DC",
X"08CA",
X"09C4",
X"09C4",
X"07D0",
X"04E2",
X"0177",
X"FD12",
X"F92A",
X"F5BF",
X"F34E",
X"F34E",
X"F542",
X"F830",
X"FC18",
X"007D",
X"04E2",
X"07D0",
X"09C4",
X"09C4",
X"08CA",
X"0659",
X"02EE",
X"FF83",
X"FC18",
X"F9A7",
X"F8AD",
X"F8AD",
X"FA24",
X"FD12",
X"00FA",
X"04E2",
X"084D",
X"0A41",
X"0ABE",
X"09C4",
X"06D6",
X"02EE",
X"FE0C",
X"F9A7",
X"F5BF",
X"F2D1",
X"F254",
X"F3CB",
X"F6B9",
X"FAA1",
X"FF83",
X"03E8",
X"0753",
X"09C4",
X"0A41",
X"0947",
X"0753",
X"03E8",
X"007D",
X"FD12",
X"FA24",
X"F830",
X"F830",
X"F92A",
X"FC18",
X"FF83",
X"03E8",
X"07D0",
X"0A41",
X"0BB8",
X"0ABE",
X"08CA",
X"04E2",
X"0000",
X"FB1E",
X"F63C",
X"F2D1",
X"F15A",
X"F254",
X"F4C5",
X"F92A",
X"FE0C",
X"0271",
X"06D6",
X"09C4",
X"0ABE",
X"0A41",
X"084D",
X"055F",
X"0177",
X"FD8F",
X"FAA1",
X"F830",
X"F736",
X"F830",
X"FAA1",
X"FE89",
X"02EE",
X"06D6",
X"0A41",
X"0BB8",
X"0C35",
X"0A41",
X"06D6",
X"0177",
X"FC18",
X"F6B9",
X"F2D1",
X"F060",
X"F0DD",
X"F34E",
X"F736",
X"FC95",
X"01F4",
X"0659",
X"09C4",
X"0BB8",
X"0BB8",
X"09C4",
X"06D6",
X"02EE",
X"FE89",
X"FB1E",
X"F830",
X"F6B9",
X"F736",
X"F92A",
X"FC95",
X"00FA",
X"055F",
X"0947",
X"0C35",
X"0D2F",
X"0C35",
X"08CA",
X"03E8",
X"FD8F",
X"F7B3",
X"F2D1",
X"EFE3",
X"EF66",
X"F15A",
X"F542",
X"FAA1",
X"007D",
X"05DC",
X"09C4",
X"0BB8",
X"0C35",
X"0ABE",
X"07D0",
X"03E8",
X"0000",
X"FB9B",
X"F8AD",
X"F6B9",
X"F63C",
X"F830",
X"FB1E",
X"FF83",
X"0465",
X"08CA",
X"0C35",
X"0DAC",
X"0DAC",
X"0B3B",
X"05DC",
X"FF83",
X"F92A",
X"F3CB",
X"EFE3",
X"EE6C",
X"EFE3",
X"F3CB",
X"F92A",
X"FF06",
X"04E2",
X"0947",
X"0BB8",
X"0CB2",
X"0BB8",
X"08CA",
X"04E2",
X"007D",
X"FC18",
X"F8AD",
X"F6B9",
X"F63C",
X"F7B3",
X"FAA1",
X"FF06",
X"036B",
X"084D",
X"0BB8",
X"0DAC",
X"0DAC",
X"0C35",
X"0753",
X"00FA",
X"FAA1",
X"F4C5",
X"F060",
X"EE6C",
X"EEE9",
X"F254",
X"F7B3",
X"FD8F",
X"036B",
X"08CA",
X"0BB8",
X"0D2F",
X"0C35",
X"09C4",
X"05DC",
X"0177",
X"FD12",
X"F92A",
X"F6B9",
X"F5BF",
X"F6B9",
X"F9A7",
X"FD8F",
X"01F4",
X"06D6",
X"0ABE",
X"0DAC",
X"0EA6",
X"0DAC",
X"09C4",
X"036B",
X"FC95",
X"F5BF",
X"F0DD",
X"ED72",
X"ED72",
X"F060",
X"F542",
X"FB9B",
X"01F4",
X"07D0",
X"0BB8",
X"0DAC",
X"0D2F",
X"0B3B",
X"0753",
X"02EE",
X"FE0C",
X"F9A7",
X"F6B9",
X"F542",
X"F5BF",
X"F830",
X"FC18",
X"00FA",
X"05DC",
X"0A41",
X"0D2F",
X"0F23",
X"0F23",
X"0BB8",
X"055F",
X"FE0C",
X"F736",
X"F1D7",
X"EDEF",
X"ECF5",
X"EEE9",
X"F3CB",
X"FA24",
X"007D",
X"06D6",
X"0ABE",
X"0D2F",
X"0DAC",
X"0BB8",
X"084D",
X"036B",
X"FF06",
X"FAA1",
X"F6B9",
X"F542",
X"F542",
X"F7B3",
X"FB1E",
X"0000",
X"055F",
X"09C4",
X"0D2F",
X"0F23",
X"0FA0",
X"0CB2",
X"06D6",
X"FF83",
X"F8AD",
X"F2D1",
X"EE6C",
X"ECF5",
X"EE6C",
X"F2D1",
X"F8AD",
X"FF83",
X"05DC",
X"0A41",
X"0D2F",
X"0DAC",
X"0CB2",
X"0947",
X"0465",
X"FF83",
X"FB1E",
X"F7B3",
X"F542",
X"F542",
X"F6B9",
X"FA24",
X"FE89",
X"03E8",
X"084D",
X"0C35",
X"0EA6",
X"101D",
X"0E29",
X"08CA",
X"0177",
X"FA24",
X"F3CB",
X"EF66",
X"ECF5",
X"ED72",
X"F15A",
X"F6B9",
X"FD8F",
X"0465",
X"09C4",
X"0CB2",
X"0E29",
X"0D2F",
X"0A41",
X"05DC",
X"00FA",
X"FC18",
X"F830",
X"F5BF",
X"F4C5",
X"F63C",
X"F92A",
X"FD12",
X"0271",
X"0753",
X"0B3B",
X"0EA6",
X"101D",
X"0F23",
X"0ABE",
X"036B",
X"FB9B",
X"F542",
X"EFE3",
X"ECF5",
X"EC78",
X"EFE3",
X"F542",
X"FC18",
X"02EE",
X"08CA",
X"0CB2",
X"0E29",
X"0DAC",
X"0B3B",
X"0753",
X"0271",
X"FD8F",
X"F8AD",
X"F5BF",
X"F448",
X"F542",
X"F7B3",
X"FB9B",
X"00FA",
X"0659",
X"0ABE",
X"0E29",
X"101D",
X"101D",
X"0C35",
X"04E2",
X"FD12",
X"F63C",
X"F0DD",
X"ECF5",
X"EBFB",
X"EE6C",
X"F3CB",
X"FA24",
X"0177",
X"07D0",
X"0C35",
X"0EA6",
X"0EA6",
X"0CB2",
X"084D",
X"036B",
X"FE89",
X"FA24",
X"F63C",
X"F448",
X"F4C5",
X"F6B9",
X"FAA1",
X"FF83",
X"04E2",
X"0947",
X"0D2F",
X"101D",
X"1117",
X"0E29",
X"07D0",
X"FF83",
X"F7B3",
X"F1D7",
X"ECF5",
X"EB7E",
X"ECF5",
X"F1D7",
X"F830",
X"FF83",
X"06D6",
X"0BB8",
X"0EA6",
X"0F23",
X"0DAC",
X"09C4",
X"0465",
X"FF83",
X"FAA1",
X"F6B9",
X"F448",
X"F448",
X"F63C",
X"F9A7",
X"FE89",
X"03E8",
X"08CA",
X"0CB2",
X"0FA0",
X"1117",
X"0F23",
X"09C4",
X"0177",
X"F92A",
X"F2D1",
X"EDEF",
X"EB01",
X"EBFB",
X"F060",
X"F6B9",
X"FE0C",
X"05DC",
X"0B3B",
X"0E29",
X"0FA0",
X"0EA6",
X"0ABE",
X"05DC",
X"007D",
X"FB9B",
X"F736",
X"F448",
X"F3CB",
X"F542",
X"F830",
X"FD12",
X"0271",
X"07D0",
X"0C35",
X"0FA0",
X"1194",
X"109A",
X"0B3B",
X"02EE",
X"FAA1",
X"F34E",
X"EDEF",
X"EA84",
X"EB7E",
X"EF66",
X"F542",
X"FD12",
X"04E2",
X"0B3B",
X"0EA6",
X"101D",
X"0F23",
X"0BB8",
X"06D6",
X"00FA",
X"FB9B",
X"F6B9",
X"F3CB",
X"F34E",
X"F4C5",
X"F7B3",
X"FC95",
X"01F4",
X"07D0",
X"0CB2",
X"101D",
X"1194",
X"1117",
X"0CB2",
X"03E8",
X"FB1E",
X"F3CB",
X"EE6C",
X"EA07",
X"EA07",
X"EDEF",
X"F448",
X"FB9B",
X"03E8",
X"0ABE",
X"0EA6",
X"109A",
X"109A",
X"0D2F",
X"084D",
X"0271",
X"FC95",
X"F736",
X"F34E",
X"F1D7",
X"F2D1",
X"F63C",
X"FB1E",
X"00FA",
X"06D6",
X"0C35",
X"101D",
X"1211",
X"1211",
X"0EA6",
X"06D6",
X"FD8F",
X"F542",
X"EEE9",
X"EA07",
X"E890",
X"EBFB",
X"F1D7",
X"F9A7",
X"01F4",
X"09C4",
X"0F23",
X"1194",
X"1194",
X"0F23",
X"0A41",
X"03E8",
X"FD8F",
X"F7B3",
X"F34E",
X"F15A",
X"F254",
X"F542",
X"FA24",
X"0000",
X"0659",
X"0BB8",
X"0FA0",
X"1211",
X"128E",
X"0FA0",
X"084D",
X"FE89",
X"F5BF",
X"EF66",
X"EA84",
X"E813",
X"EA84",
X"F0DD",
X"F830",
X"00FA",
X"0947",
X"0EA6",
X"1194",
X"1211",
X"101D",
X"0B3B",
X"04E2",
X"FE89",
X"F8AD",
X"F3CB",
X"F15A",
X"F1D7",
X"F448",
X"F92A",
X"FF06",
X"055F",
X"0B3B",
X"0FA0",
X"1211",
X"128E",
X"109A",
X"0A41",
X"007D",
X"F6B9",
X"EF66",
X"EA84",
X"E796",
X"E90D",
X"EEE9",
X"F6B9",
X"FF83",
X"084D",
X"0EA6",
X"1211",
X"130B",
X"1117",
X"0C35",
X"055F",
X"FE89",
X"F8AD",
X"F448",
X"F1D7",
X"F1D7",
X"F3CB",
X"F8AD",
X"FE89",
X"0465",
X"0A41",
X"0EA6",
X"1194",
X"1388",
X"128E",
X"0D2F",
X"02EE",
X"F830",
X"F060",
X"EA84",
X"E69C",
X"E796",
X"ED72",
X"F542",
X"FE0C",
X"0753",
X"0E29",
X"1194",
X"128E",
X"1117",
X"0CB2",
X"0659",
X"0000",
X"F9A7",
X"F542",
X"F254",
X"F1D7",
X"F34E",
X"F7B3",
X"FD12",
X"02EE",
X"08CA",
X"0DAC",
X"1194",
X"130B",
X"130B",
X"0EA6",
X"055F",
X"FAA1",
X"F1D7",
X"EB7E",
X"E796",
X"E719",
X"EBFB",
X"F34E",
X"FC18",
X"055F",
X"0D2F",
X"1117",
X"128E",
X"1194",
X"0DAC",
X"07D0",
X"00FA",
X"FAA1",
X"F5BF",
X"F254",
X"F1D7",
X"F34E",
X"F6B9",
X"FC18",
X"01F4",
X"07D0",
X"0D2F",
X"109A",
X"1211",
X"1211",
X"0FA0",
X"07D0",
X"FD12",
X"F34E",
X"ECF5",
X"E890",
X"E796",
X"EB01",
X"F254",
X"FA24",
X"02EE",
X"0B3B",
X"101D",
X"1194",
X"1117",
X"0EA6",
X"0947",
X"0271",
X"FC18",
X"F6B9",
X"F34E",
X"F254",
X"F34E",
X"F6B9",
X"FB9B",
X"00FA",
X"0659",
X"0BB8",
X"0FA0",
X"1194",
X"1211",
X"101D",
X"09C4",
X"FF06",
X"F4C5",
X"EDEF",
X"E98A",
X"E796",
X"EA84",
X"F0DD",
X"F92A",
X"01F4",
X"0A41",
X"0FA0",
X"1194",
X"1117",
X"0EA6",
X"0947",
X"02EE",
X"FD12",
X"F7B3",
X"F448",
X"F2D1",
X"F34E",
X"F63C",
X"FAA1",
X"0000",
X"055F",
X"0ABE",
X"0F23",
X"1194",
X"1211",
X"109A",
X"0B3B",
X"00FA",
X"F5BF",
X"EDEF",
X"E98A",
X"E719",
X"E90D",
X"EFE3",
X"F8AD",
X"0177",
X"09C4",
X"0FA0",
X"1211",
X"1194",
X"0F23",
X"0A41",
X"03E8",
X"FD12",
X"F830",
X"F448",
X"F254",
X"F34E",
X"F5BF",
X"FA24",
X"FF83",
X"0465",
X"0947",
X"0DAC",
X"109A",
X"1194",
X"1117",
X"0D2F",
X"03E8",
X"F8AD",
X"EF66",
X"EA84",
X"E796",
X"E813",
X"EDEF",
X"F6B9",
X"FF83",
X"084D",
X"0F23",
X"1211",
X"1194",
X"0FA0",
X"0B3B",
X"04E2",
X"FE89",
X"F92A",
X"F542",
X"F2D1",
X"F34E",
X"F4C5",
X"F8AD",
X"FE0C",
X"02EE",
X"07D0",
X"0CB2",
X"101D",
X"1211",
X"1211",
X"0FA0",
X"0753",
X"FB1E",
X"F060",
X"EA84",
X"E69C",
X"E69C",
X"EB01",
X"F3CB",
X"FD8F",
X"06D6",
X"0EA6",
X"128E",
X"128E",
X"109A",
X"0CB2",
X"0659",
X"0000",
X"F9A7",
X"F542",
X"F34E",
X"F2D1",
X"F448",
X"F7B3",
X"FC95",
X"01F4",
X"06D6",
X"0B3B",
X"0F23",
X"1194",
X"130B",
X"1194",
X"0B3B",
X"FF83",
X"F2D1",
X"EB01",
X"E719",
X"E5A2",
X"E890",
X"F15A",
X"FB1E",
X"0465",
X"0CB2",
X"1194",
X"128E",
X"1117",
X"0DAC",
X"07D0",
X"0177",
X"FB9B",
X"F6B9",
X"F448",
X"F34E",
X"F4C5",
X"F736",
X"FB1E",
X"0000",
X"04E2",
X"0947",
X"0DAC",
X"109A",
X"128E",
X"130B",
X"0EA6",
X"036B",
X"F63C",
X"ECF5",
X"E890",
X"E61F",
X"E796",
X"EEE9",
X"F8AD",
X"01F4",
X"0A41",
X"101D",
X"1211",
X"109A",
X"0DAC",
X"08CA",
X"0271",
X"FC95",
X"F830",
X"F542",
X"F448",
X"F4C5",
X"F6B9",
X"FAA1",
X"FF06",
X"036B",
X"07D0",
X"0BB8",
X"0F23",
X"109A",
X"1211",
X"109A",
X"08CA",
X"FB9B",
X"EF66",
X"E90D",
X"E69C",
X"E719",
X"EC78",
X"F542",
X"FF83",
X"08CA",
X"0F23",
X"1194",
X"1117",
X"0EA6",
X"09C4",
X"03E8",
X"FE89",
X"F92A",
X"F5BF",
X"F448",
X"F448",
X"F5BF",
X"F8AD",
X"FD8F",
X"01F4",
X"0659",
X"0ABE",
X"0EA6",
X"1117",
X"128E",
X"1194",
X"0B3B",
X"FF06",
X"F1D7",
X"EA07",
X"E69C",
X"E61F",
X"EA84",
X"F34E",
X"FD12",
X"0659",
X"0DAC",
X"1194",
X"1117",
X"0F23",
X"0B3B",
X"05DC",
X"FF83",
X"FAA1",
X"F6B9",
X"F4C5",
X"F448",
X"F542",
X"F830",
X"FC95",
X"00FA",
X"04E2",
X"0947",
X"0DAC",
X"101D",
X"1211",
X"130B",
X"0DAC",
X"0177",
X"F3CB",
X"EB7E",
X"E796",
X"E5A2",
X"E813",
X"F0DD",
X"FB1E",
X"0465",
X"0C35",
X"1117",
X"1194",
X"101D",
X"0CB2",
X"06D6",
X"00FA",
X"FB1E",
X"F736",
X"F542",
X"F4C5",
X"F5BF",
X"F7B3",
X"FC18",
X"007D",
X"04E2",
X"08CA",
X"0C35",
X"0EA6",
X"109A",
X"1211",
X"0FA0",
X"05DC",
X"F7B3",
X"EC78",
X"E796",
X"E69C",
X"E813",
X"EEE9",
X"F8AD",
X"0271",
X"0ABE",
X"101D",
X"1194",
X"101D",
X"0D2F",
X"07D0",
X"0177",
X"FB9B",
X"F7B3",
X"F5BF",
X"F542",
X"F5BF",
X"F7B3",
X"FB1E",
X"FF83",
X"036B",
X"0753",
X"0ABE",
X"0E29",
X"101D",
X"1211",
X"1194",
X"09C4",
X"FC95",
X"EFE3",
X"E890",
X"E61F",
X"E69C",
X"EB7E",
X"F4C5",
X"FF06",
X"084D",
X"0FA0",
X"128E",
X"1194",
X"0EA6",
X"09C4",
X"036B",
X"FD12",
X"F830",
X"F5BF",
X"F542",
X"F5BF",
X"F7B3",
X"FAA1",
X"FE89",
X"01F4",
X"055F",
X"08CA",
X"0CB2",
X"0FA0",
X"128E",
X"1388",
X"0E29",
X"00FA",
X"F2D1",
X"EA07",
X"E61F",
X"E525",
X"E890",
X"F15A",
X"FB9B",
X"055F",
X"0DAC",
X"128E",
X"128E",
X"109A",
X"0BB8",
X"05DC",
X"FF06",
X"F92A",
X"F5BF",
X"F448",
X"F4C5",
X"F6B9",
X"F9A7",
X"FD12",
X"00FA",
X"04E2",
X"07D0",
X"0BB8",
X"0F23",
X"1194",
X"1405",
X"1117",
X"05DC",
X"F6B9",
X"EB01",
X"E61F",
X"E4A8",
X"E69C",
X"EDEF",
X"F92A",
X"036B",
X"0C35",
X"128E",
X"1388",
X"1194",
X"0DAC",
X"07D0",
X"007D",
X"F9A7",
X"F63C",
X"F4C5",
X"F4C5",
X"F5BF",
X"F8AD",
X"FC95",
X"007D",
X"036B",
X"06D6",
X"0ABE",
X"0E29",
X"109A",
X"130B",
X"128E",
X"0A41",
X"FB1E",
X"ED72",
X"E719",
X"E4A8",
X"E525",
X"EB01",
X"F5BF",
X"007D",
X"0A41",
X"1194",
X"1482",
X"128E",
X"0F23",
X"09C4",
X"0271",
X"FB1E",
X"F6B9",
X"F4C5",
X"F448",
X"F542",
X"F7B3",
X"FB1E",
X"FF83",
X"02EE",
X"05DC",
X"0947",
X"0D2F",
X"0F23",
X"1117",
X"130B",
X"0EA6",
X"01F4",
X"F2D1",
X"E90D",
X"E525",
X"E4A8",
X"E813",
X"F15A",
X"FC95",
X"06D6",
X"0FA0",
X"1482",
X"1388",
X"0FA0",
X"0ABE",
X"0465",
X"FD8F",
X"F830",
X"F542",
X"F448",
X"F542",
X"F736",
X"F9A7",
X"FD12",
X"00FA",
X"0465",
X"0753",
X"0ABE",
X"0E29",
X"109A",
X"1388",
X"1388",
X"0A41",
X"F9A7",
X"EBFB",
X"E5A2",
X"E42B",
X"E525",
X"EB01",
X"F6B9",
X"0271",
X"0C35",
X"130B",
X"1482",
X"1211",
X"0DAC",
X"084D",
X"007D",
X"F9A7",
X"F5BF",
X"F3CB",
X"F448",
X"F6B9",
X"F8AD",
X"FB9B",
X"FF83",
X"02EE",
X"0659",
X"09C4",
X"0D2F",
X"0FA0",
X"130B",
X"15F9",
X"109A",
X"0177",
X"EFE3",
X"E61F",
X"E331",
X"E331",
X"E69C",
X"F0DD",
X"FD8F",
X"08CA",
X"1117",
X"157C",
X"1405",
X"101D",
X"0ABE",
X"036B",
X"FC95",
X"F7B3",
X"F4C5",
X"F3CB",
X"F542",
X"F736",
X"FAA1",
X"FE0C",
X"0177",
X"03E8",
X"0753",
X"0BB8",
X"0F23",
X"1194",
X"14FF",
X"1405",
X"0947",
X"F7B3",
X"E98A",
X"E331",
X"E237",
X"E4A8",
X"EBFB",
X"F830",
X"0465",
X"0DAC",
X"1405",
X"14FF",
X"1211",
X"0E29",
X"0753",
X"FF06",
X"F92A",
X"F542",
X"F3CB",
X"F3CB",
X"F5BF",
X"F830",
X"FC18",
X"FF83",
X"0271",
X"055F",
X"0947",
X"0E29",
X"1194",
X"14FF",
X"17ED",
X"1211",
X"00FA",
X"EE6C",
X"E42B",
X"E13D",
X"E237",
X"E69C",
X"F15A",
X"FF06",
X"0A41",
X"128E",
X"1676",
X"1482",
X"0FA0",
X"0A41",
X"0271",
X"FB1E",
X"F6B9",
X"F448",
X"F34E",
X"F448",
X"F6B9",
X"FAA1",
X"FE89",
X"0271",
X"055F",
X"08CA",
X"0CB2",
X"101D",
X"130B",
X"15F9",
X"1388",
X"0659",
X"F4C5",
X"E796",
X"E2B4",
X"E237",
X"E525",
X"EE6C",
X"FB9B",
X"06D6",
X"0F23",
X"157C",
X"15F9",
X"1211",
X"0CB2",
X"04E2",
X"FC95",
X"F6B9",
X"F448",
X"F34E",
X"F3CB",
X"F5BF",
X"F92A",
X"FD8F",
X"0177",
X"0465",
X"0753",
X"0A41",
X"0E29",
X"1117",
X"1388",
X"1388",
X"0BB8",
X"FD12",
X"EDEF",
X"E5A2",
X"E237",
X"E3AE",
X"E98A",
X"F542",
X"01F4",
X"0BB8",
X"1388",
X"16F3",
X"14FF",
X"0FA0",
X"08CA",
X"007D",
X"F9A7",
X"F5BF",
X"F3CB",
X"F34E",
X"F3CB",
X"F6B9",
X"FA24",
X"FE0C",
X"0177",
X"04E2",
X"0947",
X"0DAC",
X"1117",
X"1388",
X"15F9",
X"130B",
X"06D6",
X"F5BF",
X"E813",
X"E1BA",
X"E0C0",
X"E4A8",
X"ED72",
X"FAA1",
X"0659",
X"0FA0",
X"15F9",
X"1676",
X"1194",
X"0C35",
X"055F",
X"FD8F",
X"F7B3",
X"F4C5",
X"F3CB",
X"F3CB",
X"F5BF",
X"F8AD",
X"FC18",
X"FF06",
X"01F4",
X"05DC",
X"09C4",
X"0DAC",
X"1194",
X"14FF",
X"186A",
X"128E",
X"0271",
X"F060",
X"E4A8",
X"E043",
X"E13D",
X"E69C",
X"F15A",
X"FF83",
X"0B3B",
X"130B",
X"1770",
X"157C",
X"0F23",
X"08CA",
X"007D",
X"F9A7",
X"F5BF",
X"F4C5",
X"F448",
X"F542",
X"F7B3",
X"FB1E",
X"FD8F",
X"FF83",
X"0271",
X"055F",
X"09C4",
X"0E29",
X"1211",
X"1770",
X"1964",
X"101D",
X"FD12",
X"EA84",
X"E13D",
X"DF49",
X"E1BA",
X"E90D",
X"F63C",
X"04E2",
X"0F23",
X"15F9",
X"17ED",
X"1405",
X"0D2F",
X"04E2",
X"FC95",
X"F6B9",
X"F4C5",
X"F4C5",
X"F5BF",
X"F7B3",
X"FA24",
X"FC18",
X"FE0C",
X"FF83",
X"0271",
X"0659",
X"0B3B",
X"101D",
X"14FF",
X"1A5E",
X"16F3",
X"07D0",
X"F3CB",
X"E42B",
X"DE4F",
X"DECC",
X"E42B",
X"EEE9",
X"FD8F",
X"0ABE",
X"1388",
X"186A",
X"16F3",
X"101D",
X"08CA",
X"007D",
X"F92A",
X"F542",
X"F3CB",
X"F4C5",
X"F5BF",
X"F7B3",
X"FAA1",
X"FD8F",
X"FF06",
X"0177",
X"055F",
X"0ABE",
X"0FA0",
X"1388",
X"18E7",
X"1ADB",
X"101D",
X"FB9B",
X"E890",
X"DECC",
X"DDD2",
X"E13D",
X"E98A",
X"F6B9",
X"05DC",
X"109A",
X"16F3",
X"186A",
X"1388",
X"0C35",
X"0465",
X"FC95",
X"F6B9",
X"F4C5",
X"F5BF",
X"F6B9",
X"F7B3",
X"F92A",
X"FB9B",
X"FE0C",
X"FF83",
X"01F4",
X"05DC",
X"0B3B",
X"101D",
X"14FF",
X"19E1",
X"1770",
X"08CA",
X"F542",
X"E5A2",
X"DECC",
X"DECC",
X"E3AE",
X"EDEF",
X"FC95",
X"09C4",
X"128E",
X"1770",
X"16F3",
X"1117",
X"09C4",
X"00FA",
X"F92A",
X"F5BF",
X"F542",
X"F63C",
X"F736",
X"F8AD",
X"FAA1",
X"FC95",
X"FE89",
X"0000",
X"036B",
X"0753",
X"0C35",
X"109A",
X"15F9",
X"1A5E",
X"1482",
X"03E8",
X"EFE3",
X"E2B4",
X"DECC",
X"DFC6",
X"E61F",
X"F1D7",
X"00FA",
X"0D2F",
X"157C",
X"186A",
X"14FF",
X"0E29",
X"0659",
X"FE0C",
X"F7B3",
X"F4C5",
X"F4C5",
X"F6B9",
X"F8AD",
X"FAA1",
X"FC95",
X"FE0C",
X"FF06",
X"007D",
X"03E8",
X"08CA",
X"0DAC",
X"1211",
X"17ED",
X"1964",
X"0E29",
X"FA24",
X"E813",
X"DFC6",
X"DF49",
X"E331",
X"EB7E",
X"FA24",
X"084D",
X"1211",
X"1770",
X"1676",
X"1117",
X"09C4",
X"01F4",
X"FA24",
X"F5BF",
X"F448",
X"F4C5",
X"F6B9",
X"F92A",
X"FB1E",
X"FD8F",
X"FF06",
X"007D",
X"03E8",
X"084D",
X"0CB2",
X"1117",
X"1676",
X"1ADB",
X"1482",
X"0271",
X"ECF5",
X"E043",
X"DDD2",
X"E0C0",
X"E796",
X"F34E",
X"0271",
X"0E29",
X"157C",
X"17ED",
X"1482",
X"0DAC",
X"0659",
X"FE0C",
X"F736",
X"F448",
X"F448",
X"F63C",
X"F7B3",
X"FA24",
X"FC18",
X"FE89",
X"007D",
X"01F4",
X"04E2",
X"08CA",
X"0DAC",
X"1211",
X"17ED",
X"186A",
X"0CB2",
X"FA24",
X"E90D",
X"E043",
X"DF49",
X"E2B4",
X"EBFB",
X"F9A7",
X"0753",
X"109A",
X"1676",
X"16F3",
X"1211",
X"0B3B",
X"036B",
X"FB1E",
X"F63C",
X"F4C5",
X"F542",
X"F736",
X"F8AD",
X"FA24",
X"FC18",
X"FD8F",
X"FF83",
X"02EE",
X"06D6",
X"0ABE",
X"0EA6",
X"1388",
X"18E7",
X"18E7",
X"0BB8",
X"F7B3",
X"E61F",
X"DECC",
X"DECC",
X"E3AE",
X"ED72",
X"FB1E",
X"084D",
X"128E",
X"16F3",
X"15F9",
X"101D",
X"08CA",
X"00FA",
X"FA24",
X"F63C",
X"F5BF",
X"F63C",
X"F7B3",
X"F92A",
X"FB9B",
X"FC95",
X"FD12",
X"FF06",
X"02EE",
X"0753",
X"0C35",
X"109A",
X"1676",
X"1C52",
X"18E7",
X"0753",
X"F0DD",
X"E13D",
X"DD55",
X"DF49",
X"E5A2",
X"F0DD",
X"0000",
X"0D2F",
X"1482",
X"1676",
X"1405",
X"0D2F",
X"055F",
X"FE0C",
X"F8AD",
X"F63C",
X"F63C",
X"F7B3",
X"F9A7",
X"FAA1",
X"FC18",
X"FC95",
X"FD8F",
X"FF83",
X"02EE",
X"06D6",
X"0ABE",
X"0EA6",
X"1482",
X"1BD5",
X"1ADB",
X"0947",
X"F15A",
X"DFC6",
X"DB61",
X"DECC",
X"E61F",
X"F15A",
X"00FA",
X"0EA6",
X"157C",
X"1770",
X"1482",
X"0C35",
X"02EE",
X"FC18",
X"F7B3",
X"F6B9",
X"F7B3",
X"F9A7",
X"FB1E",
X"FC95",
X"FC18",
X"FB1E",
X"FB1E",
X"FD12",
X"00FA",
X"05DC",
X"0B3B",
X"109A",
X"17ED",
X"2134",
X"1DC9",
X"06D6",
X"EB7E",
X"DB61",
X"D96D",
X"DE4F",
X"E69C",
X"F1D7",
X"036B",
X"1211",
X"1770",
X"17ED",
X"1405",
X"0ABE",
X"00FA",
X"FAA1",
X"F63C",
X"F542",
X"F6B9",
X"FA24",
X"FC95",
X"FD8F",
X"FC95",
X"FC18",
X"FC95",
X"FE89",
X"0271",
X"06D6",
X"0C35",
X"1117",
X"17ED",
X"20B7",
X"1A5E",
X"0271",
X"E813",
X"DA67",
X"DA67",
X"E043",
X"E890",
X"F542",
X"06D6",
X"14FF",
X"18E7",
X"1676",
X"1117",
X"084D",
X"FF83",
X"F8AD",
X"F448",
X"F4C5",
X"F830",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"007D",
X"0465",
X"084D",
X"0CB2",
X"109A",
X"17ED",
X"1FBD",
X"1770",
X"FE0C",
X"E525",
X"D96D",
X"DA67",
X"E0C0",
X"EA07",
X"F7B3",
X"0ABE",
X"16F3",
X"19E1",
X"16F3",
X"109A",
X"0753",
X"FE0C",
X"F6B9",
X"F34E",
X"F448",
X"F830",
X"FB1E",
X"FB9B",
X"FB1E",
X"FC18",
X"FD8F",
X"FE89",
X"00FA",
X"04E2",
X"0947",
X"0DAC",
X"1117",
X"1770",
X"2134",
X"1964",
X"FF83",
X"E525",
X"D873",
X"D9EA",
X"E043",
X"E90D",
X"F6B9",
X"0ABE",
X"186A",
X"1A5E",
X"1676",
X"0FA0",
X"06D6",
X"FD8F",
X"F6B9",
X"F34E",
X"F4C5",
X"F830",
X"FB1E",
X"FB1E",
X"FB9B",
X"FC95",
X"FC95",
X"FD8F",
X"007D",
X"04E2",
X"0947",
X"0DAC",
X"101D",
X"14FF",
X"203A",
X"1CCF",
X"036B",
X"E796",
X"D7F6",
X"D873",
X"E0C0",
X"E98A",
X"F5BF",
X"0947",
X"18E7",
X"1A5E",
X"15F9",
X"0F23",
X"0659",
X"FD12",
X"F5BF",
X"F34E",
X"F542",
X"F92A",
X"FB1E",
X"FB9B",
X"FC18",
X"FD12",
X"FD12",
X"FD8F",
X"0000",
X"0465",
X"084D",
X"0CB2",
X"101D",
X"1405",
X"1FBD",
X"1FBD",
X"084D",
X"EA84",
X"D7F6",
X"D67F",
X"DE4F",
X"E890",
X"F3CB",
X"06D6",
X"17ED",
X"1BD5",
X"16F3",
X"0FA0",
X"0659",
X"FD12",
X"F63C",
X"F3CB",
X"F4C5",
X"F830",
X"FB1E",
X"FB9B",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"0000",
X"0465",
X"09C4",
X"0E29",
X"1117",
X"130B",
X"1E46",
X"203A",
X"0B3B",
X"ED72",
X"D873",
X"D585",
X"DC5B",
X"E796",
X"F3CB",
X"05DC",
X"16F3",
X"1B58",
X"1676",
X"0F23",
X"06D6",
X"FD12",
X"F5BF",
X"F3CB",
X"F63C",
X"F9A7",
X"FB9B",
X"FB1E",
X"FA24",
X"FB9B",
X"FC95",
X"FD12",
X"0000",
X"0465",
X"0947",
X"0CB2",
X"0FA0",
X"128E",
X"1DC9",
X"23A5",
X"0FA0",
X"F060",
X"D8F0",
X"D40E",
X"DBDE",
X"E719",
X"F1D7",
X"01F4",
X"1482",
X"1BD5",
X"17ED",
X"101D",
X"0753",
X"FC95",
X"F5BF",
X"F3CB",
X"F6B9",
X"FB1E",
X"FC95",
X"FB9B",
X"FAA1",
X"FB9B",
X"FC95",
X"FC95",
X"FE89",
X"0271",
X"084D",
X"0C35",
X"0F23",
X"109A",
X"19E1",
X"22AB",
X"130B",
X"F5BF",
X"DD55",
X"D67F",
X"DC5B",
X"E796",
X"F1D7",
X"0000",
X"1211",
X"19E1",
X"17ED",
X"101D",
X"0753",
X"FD12",
X"F5BF",
X"F34E",
X"F5BF",
X"FA24",
X"FC95",
X"FE0C",
X"FC95",
X"FD8F",
X"FE89",
X"FD8F",
X"FE89",
X"00FA",
X"055F",
X"0947",
X"0CB2",
X"0EA6",
X"15F9",
X"21B1",
X"17ED",
X"FD12",
X"E331",
X"D7F6",
X"DBDE",
X"E5A2",
X"F0DD",
X"FC95",
X"0DAC",
X"186A",
X"17ED",
X"1117",
X"08CA",
X"FF83",
X"F6B9",
X"F34E",
X"F448",
X"F92A",
X"FC18",
X"FD8F",
X"FD8F",
X"FE0C",
X"FF06",
X"FE89",
X"FF83",
X"0177",
X"055F",
X"08CA",
X"0B3B",
X"0CB2",
X"0FA0",
X"1C52",
X"1D4C",
X"08CA",
X"ECF5",
X"DB61",
X"DA67",
X"E237",
X"EDEF",
X"F830",
X"0659",
X"1482",
X"1770",
X"128E",
X"0BB8",
X"02EE",
X"F9A7",
X"F4C5",
X"F448",
X"F736",
X"FAA1",
X"FC18",
X"FD12",
X"FD8F",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"03E8",
X"084D",
X"0BB8",
X"0D2F",
X"0F23",
X"18E7",
X"1FBD",
X"0F23",
X"F2D1",
X"DDD2",
X"D8F0",
X"DFC6",
X"EB01",
X"F5BF",
X"036B",
X"1194",
X"17ED",
X"1405",
X"0D2F",
X"04E2",
X"FB1E",
X"F448",
X"F34E",
X"F5BF",
X"F9A7",
X"FB1E",
X"FC18",
X"FD12",
X"FE89",
X"FF06",
X"FF06",
X"00FA",
X"0465",
X"084D",
X"0A41",
X"0C35",
X"0EA6",
X"19E1",
X"222E",
X"1117",
X"F448",
X"DCD8",
X"D779",
X"DDD2",
X"E890",
X"F448",
X"0271",
X"130B",
X"1964",
X"1676",
X"0F23",
X"05DC",
X"FB9B",
X"F4C5",
X"F254",
X"F4C5",
X"F92A",
X"FB9B",
X"FC95",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"00FA",
X"036B",
X"084D",
X"0BB8",
X"0D2F",
X"0FA0",
X"18E7",
X"21B1",
X"1194",
X"F3CB",
X"DC5B",
X"D585",
X"DCD8",
X"E890",
X"F448",
X"0271",
X"1388",
X"1B58",
X"17ED",
X"101D",
X"0659",
X"FB9B",
X"F448",
X"F2D1",
X"F3CB",
X"F736",
X"FAA1",
X"FC95",
X"FD8F",
X"FE89",
X"FF83",
X"FE89",
X"007D",
X"02EE",
X"0659",
X"0947",
X"0C35",
X"0EA6",
X"186A",
X"2422",
X"17ED",
X"FB9B",
X"E043",
X"D585",
X"D96D",
X"E42B",
X"F060",
X"FE0C",
X"1117",
X"1BD5",
X"1964",
X"1117",
X"0753",
X"FD8F",
X"F4C5",
X"F15A",
X"F34E",
X"F736",
X"FB1E",
X"FD12",
X"FD8F",
X"FF83",
X"007D",
X"FE89",
X"FF06",
X"01F4",
X"04E2",
X"0753",
X"0B3B",
X"0E29",
X"1388",
X"203A",
X"1EC3",
X"07D0",
X"EB7E",
X"D8F0",
X"D67F",
X"DFC6",
X"ECF5",
X"F9A7",
X"09C4",
X"18E7",
X"1B58",
X"1388",
X"09C4",
X"0000",
X"F7B3",
X"F2D1",
X"F34E",
X"F63C",
X"F9A7",
X"FC18",
X"FD12",
X"FF06",
X"01F4",
X"0000",
X"FE0C",
X"FE89",
X"007D",
X"0465",
X"07D0",
X"0C35",
X"0FA0",
X"1A5E",
X"2422",
X"157C",
X"F8AD",
X"DF49",
X"D602",
X"DB61",
X"E813",
X"F4C5",
X"02EE",
X"1388",
X"1ADB",
X"157C",
X"0B3B",
X"0271",
X"F9A7",
X"F448",
X"F3CB",
X"F63C",
X"FAA1",
X"FE0C",
X"FF83",
X"0000",
X"00FA",
X"0000",
X"FD12",
X"FD12",
X"FE0C",
X"02EE",
X"0753",
X"0B3B",
X"0E29",
X"15F9",
X"2328",
X"1C52",
X"01F4",
X"E61F",
X"D67F",
X"D7F6",
X"E42B",
X"F0DD",
X"FD12",
X"0DAC",
X"1964",
X"186A",
X"0F23",
X"05DC",
X"FC18",
X"F542",
X"F448",
X"F7B3",
X"FC18",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"FD8F",
X"FC95",
X"FC95",
X"FE89",
X"036B",
X"07D0",
X"0C35",
X"1117",
X"1F40",
X"222E",
X"0C35",
X"EF66",
X"D9EA",
X"D779",
X"E0C0",
X"EE6C",
X"FA24",
X"06D6",
X"1388",
X"1770",
X"109A",
X"06D6",
X"FE0C",
X"F736",
X"F448",
X"F6B9",
X"FB9B",
X"FE89",
X"FF83",
X"007D",
X"0271",
X"01F4",
X"FD12",
X"FAA1",
X"FC18",
X"FE89",
X"03E8",
X"08CA",
X"0BB8",
X"0E29",
X"16F3",
X"20B7",
X"1676",
X"FD12",
X"E331",
X"D873",
X"DD55",
X"E90D",
X"F542",
X"00FA",
X"0EA6",
X"15F9",
X"1211",
X"08CA",
X"007D",
X"F92A",
X"F5BF",
X"F63C",
X"F9A7",
X"FE89",
X"007D",
X"007D",
X"0177",
X"01F4",
X"0000",
X"FB9B",
X"FAA1",
X"FC95",
X"007D",
X"0659",
X"0A41",
X"0CB2",
X"1117",
X"1D4C",
X"21B1",
X"0EA6",
X"F254",
X"DDD2",
X"D9EA",
X"E1BA",
X"EE6C",
X"F9A7",
X"055F",
X"1194",
X"130B",
X"0B3B",
X"0271",
X"FB9B",
X"F6B9",
X"F63C",
X"F8AD",
X"FC95",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"00FA",
X"FE0C",
X"FA24",
X"FAA1",
X"FE0C",
X"03E8",
X"08CA",
X"0BB8",
X"0E29",
X"157C",
X"2328",
X"1D4C",
X"0271",
X"E719",
X"D96D",
X"DB61",
X"E5A2",
X"F448",
X"FF06",
X"0B3B",
X"130B",
X"0EA6",
X"055F",
X"FE0C",
X"FA24",
X"F7B3",
X"F7B3",
X"FAA1",
X"FE89",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"FF06",
X"FC18",
X"FB1E",
X"FC95",
X"00FA",
X"0659",
X"09C4",
X"0C35",
X"0EA6",
X"1964",
X"222E",
X"14FF",
X"F92A",
X"E331",
X"DB61",
X"DFC6",
X"EB7E",
X"F736",
X"00FA",
X"0C35",
X"1194",
X"0B3B",
X"01F4",
X"FC95",
X"FA24",
X"F9A7",
X"FA24",
X"FD12",
X"0000",
X"00FA",
X"00FA",
X"0000",
X"FE89",
X"FD12",
X"FB1E",
X"FB1E",
X"FE89",
X"02EE",
X"0753",
X"09C4",
X"0C35",
X"1117",
X"1DC9",
X"23A5",
X"109A",
X"F448",
X"E0C0",
X"DC5B",
X"E331",
X"EEE9",
X"F830",
X"00FA",
X"0C35",
X"0EA6",
X"0753",
X"0000",
X"FD8F",
X"FC18",
X"FAA1",
X"FC18",
X"FF83",
X"0177",
X"00FA",
X"0000",
X"FE89",
X"FE0C",
X"FC18",
X"F92A",
X"FAA1",
X"FF83",
X"04E2",
X"084D",
X"0A41",
X"0DAC",
X"1388",
X"1F40",
X"2134",
X"0BB8",
X"F0DD",
X"DFC6",
X"DDD2",
X"E5A2",
X"EF66",
X"F7B3",
X"00FA",
X"0ABE",
X"0B3B",
X"03E8",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FE89",
X"0177",
X"02EE",
X"0177",
X"FF06",
X"FD8F",
X"FC95",
X"FAA1",
X"F9A7",
X"FC95",
X"01F4",
X"0659",
X"0947",
X"0ABE",
X"0DAC",
X"157C",
X"22AB",
X"1E46",
X"0465",
X"EB01",
X"DDD2",
X"DECC",
X"E719",
X"F060",
X"F830",
X"01F4",
X"0B3B",
X"09C4",
X"02EE",
X"007D",
X"00FA",
X"FF83",
X"FE0C",
X"0000",
X"01F4",
X"0177",
X"FF06",
X"FD12",
X"FB9B",
X"FAA1",
X"FA24",
X"FB1E",
X"0000",
X"05DC",
X"07D0",
X"08CA",
X"0ABE",
X"0DAC",
X"18E7",
X"2710",
X"1B58",
X"FD8F",
X"E525",
X"DAE4",
X"DE4F",
X"E796",
X"F1D7",
X"F8AD",
X"0465",
X"0C35",
X"07D0",
X"01F4",
X"00FA",
X"0271",
X"0000",
X"FF06",
X"007D",
X"0271",
X"00FA",
X"FD8F",
X"FB1E",
X"FAA1",
X"FB9B",
X"FA24",
X"FC18",
X"01F4",
X"06D6",
X"0947",
X"0A41",
X"0CB2",
X"109A",
X"1FBD",
X"2616",
X"101D",
X"F2D1",
X"DF49",
X"DBDE",
X"E0C0",
X"EA84",
X"F2D1",
X"FB9B",
X"084D",
X"0BB8",
X"05DC",
X"01F4",
X"0271",
X"0271",
X"007D",
X"007D",
X"01F4",
X"0177",
X"FE0C",
X"FB1E",
X"FAA1",
X"FC95",
X"FC95",
X"FB1E",
X"FE89",
X"04E2",
X"08CA",
X"08CA",
X"084D",
X"0A41",
X"101D",
X"1DC9",
X"22AB",
X"0E29",
X"F254",
X"E0C0",
X"DC5B",
X"E13D",
X"EB01",
X"F4C5",
X"FE0C",
X"0947",
X"0C35",
X"05DC",
X"01F4",
X"0271",
X"01F4",
X"FF83",
X"FF06",
X"007D",
X"FF83",
X"FC18",
X"FB1E",
X"FB9B",
X"FD8F",
X"FE0C",
X"FD12",
X"0000",
X"03E8",
X"05DC",
X"06D6",
X"07D0",
X"0B3B",
X"109A",
X"1E46",
X"22AB",
X"0EA6",
X"F34E",
X"E0C0",
X"DB61",
X"E13D",
X"EBFB",
X"F542",
X"FE89",
X"07D0",
X"0947",
X"04E2",
X"02EE",
X"03E8",
X"01F4",
X"FF06",
X"FE0C",
X"0000",
X"FF83",
X"FC18",
X"FB9B",
X"FD12",
X"FF83",
X"FF06",
X"FE0C",
X"007D",
X"04E2",
X"0753",
X"06D6",
X"0659",
X"0A41",
X"128E",
X"203A",
X"21B1",
X"0A41",
X"EF66",
X"DF49",
X"DB61",
X"E237",
X"EC78",
X"F6B9",
X"00FA",
X"0A41",
X"09C4",
X"04E2",
X"036B",
X"0465",
X"01F4",
X"FE89",
X"FE0C",
X"FF06",
X"FE0C",
X"FB9B",
X"FB9B",
X"FD8F",
X"FF83",
X"FF83",
X"FE89",
X"0271",
X"055F",
X"05DC",
X"055F",
X"0659",
X"0A41",
X"1194",
X"1F40",
X"203A",
X"08CA",
X"EF66",
X"DE4F",
X"DB61",
X"E331",
X"EE6C",
X"F7B3",
X"00FA",
X"09C4",
X"0ABE",
X"0753",
X"055F",
X"0465",
X"0000",
X"FC95",
X"FD12",
X"FE0C",
X"FD12",
X"FC95",
X"FE89",
X"0000",
X"0000",
X"FE89",
X"FC95",
X"007D",
X"03E8",
X"0465",
X"04E2",
X"0659",
X"0ABE",
X"1388",
X"222E",
X"203A",
X"0659",
X"EC78",
X"DC5B",
X"DAE4",
X"E3AE",
X"EEE9",
X"F8AD",
X"02EE",
X"0BB8",
X"0B3B",
X"0753",
X"055F",
X"0465",
X"FF06",
X"FB9B",
X"FC95",
X"FD8F",
X"FC95",
X"FD12",
X"0000",
X"0177",
X"01F4",
X"FF06",
X"FC18",
X"0000",
X"0271",
X"02EE",
X"0465",
X"07D0",
X"0C35",
X"1770",
X"251C",
X"1B58",
X"FF83",
X"E796",
X"DAE4",
X"DCD8",
X"E69C",
X"F0DD",
X"F9A7",
X"055F",
X"0D2F",
X"0ABE",
X"0659",
X"055F",
X"03E8",
X"FF83",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FE89",
X"0177",
X"01F4",
X"007D",
X"FC95",
X"FC18",
X"0000",
X"01F4",
X"02EE",
X"0465",
X"084D",
X"0FA0",
X"1CCF",
X"2422",
X"1211",
X"F6B9",
X"E331",
X"DC5B",
X"E0C0",
X"EA84",
X"F3CB",
X"FD8F",
X"0947",
X"0D2F",
X"084D",
X"055F",
X"055F",
X"0271",
X"FD8F",
X"FB1E",
X"FD12",
X"FE0C",
X"FD12",
X"FD8F",
X"FF06",
X"00FA",
X"007D",
X"FD8F",
X"FE89",
X"0271",
X"0465",
X"03E8",
X"04E2",
X"08CA",
X"109A",
X"1FBD",
X"20B7",
X"08CA",
X"EEE9",
X"DECC",
X"DB61",
X"E331",
X"EE6C",
X"F7B3",
X"0271",
X"0DAC",
X"0DAC",
X"08CA",
X"05DC",
X"03E8",
X"0000",
X"FC18",
X"FB1E",
X"FD12",
X"FD8F",
X"FC18",
X"FD12",
X"0000",
X"0177",
X"007D",
X"FE89",
X"007D",
X"03E8",
X"055F",
X"04E2",
X"05DC",
X"09C4",
X"1117",
X"1E46",
X"1C52",
X"0465",
X"EBFB",
X"DDD2",
X"DCD8",
X"E525",
X"EFE3",
X"F8AD",
X"036B",
X"0D2F",
X"0D2F",
X"07D0",
X"04E2",
X"036B",
X"FF83",
X"FD12",
X"FC18",
X"FD12",
X"FD8F",
X"FD12",
X"FE89",
X"0000",
X"00FA",
X"0000",
X"FF06",
X"0177",
X"02EE",
X"0465",
X"055F",
X"0753",
X"0A41",
X"130B",
X"1F40",
X"1A5E",
X"01F4",
X"EA07",
X"DDD2",
X"DE4F",
X"E719",
X"F15A",
X"FAA1",
X"05DC",
X"0DAC",
X"0C35",
X"07D0",
X"04E2",
X"0271",
X"FE89",
X"FAA1",
X"FAA1",
X"FC18",
X"FB9B",
X"FC18",
X"FF83",
X"0177",
X"01F4",
X"00FA",
X"007D",
X"0177",
X"02EE",
X"036B",
X"0465",
X"05DC",
X"0B3B",
X"16F3",
X"2134",
X"157C",
X"FC18",
X"E69C",
X"DD55",
X"E043",
X"E90D",
X"F2D1",
X"FC18",
X"08CA",
X"0E29",
X"09C4",
X"05DC",
X"03E8",
X"01F4",
X"FE0C",
X"FB9B",
X"FC95",
X"FD8F",
X"FD12",
X"FE0C",
X"00FA",
X"0271",
X"0177",
X"FF83",
X"FF06",
X"00FA",
X"0271",
X"0271",
X"02EE",
X"06D6",
X"0F23",
X"1C52",
X"1EC3",
X"0B3B",
X"F2D1",
X"E237",
X"DF49",
X"E525",
X"ECF5",
X"F4C5",
X"FF06",
X"0B3B",
X"0D2F",
X"08CA",
X"05DC",
X"03E8",
X"0177",
X"FE0C",
X"FC95",
X"FD8F",
X"FD8F",
X"FD12",
X"FF06",
X"01F4",
X"02EE",
X"00FA",
X"FE89",
X"FF06",
X"01F4",
X"0271",
X"0177",
X"036B",
X"08CA",
X"15F9",
X"2328",
X"18E7",
X"0000",
X"EA07",
X"DECC",
X"E13D",
X"E890",
X"EF66",
X"F7B3",
X"04E2",
X"0D2F",
X"0ABE",
X"06D6",
X"0465",
X"02EE",
X"00FA",
X"FE0C",
X"FD8F",
X"FE0C",
X"FD12",
X"FC18",
X"FE89",
X"00FA",
X"0177",
X"FF83",
X"FF83",
X"01F4",
X"0465",
X"0465",
X"03E8",
X"05DC",
X"0D2F",
X"1D4C",
X"222E",
X"0D2F",
X"F3CB",
X"E1BA",
X"DDD2",
X"E3AE",
X"EB7E",
X"F34E",
X"FD8F",
X"0ABE",
X"0EA6",
X"09C4",
X"055F",
X"036B",
X"0177",
X"FF06",
X"FD12",
X"FD8F",
X"FD8F",
X"FB9B",
X"FC95",
X"FF06",
X"0177",
X"00FA",
X"FF83",
X"007D",
X"036B",
X"055F",
X"0465",
X"0465",
X"0753",
X"1194",
X"1F40",
X"1ADB",
X"036B",
X"ECF5",
X"E043",
X"E0C0",
X"E796",
X"EEE9",
X"F6B9",
X"02EE",
X"0DAC",
X"0CB2",
X"0753",
X"0465",
X"0271",
X"007D",
X"FE89",
X"FD8F",
X"FE0C",
X"FD8F",
X"FC18",
X"FD12",
X"0000",
X"0177",
X"0000",
X"FE89",
X"007D",
X"02EE",
X"03E8",
X"036B",
X"03E8",
X"0A41",
X"1770",
X"21B1",
X"1770",
X"FE0C",
X"E890",
X"DF49",
X"E237",
X"E98A",
X"F0DD",
X"FAA1",
X"0753",
X"0F23",
X"0B3B",
X"05DC",
X"02EE",
X"0177",
X"0000",
X"FD8F",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FF06",
X"01F4",
X"0177",
X"FF06",
X"FE89",
X"007D",
X"02EE",
X"02EE",
X"036B",
X"0753",
X"1117",
X"1EC3",
X"1FBD",
X"0B3B",
X"F1D7",
X"E0C0",
X"DE4F",
X"E5A2",
X"EEE9",
X"F6B9",
X"007D",
X"0CB2",
X"0EA6",
X"09C4",
X"055F",
X"0177",
X"FF06",
X"FE0C",
X"FD8F",
X"FC18",
X"FC18",
X"FB9B",
X"FC95",
X"007D",
X"02EE",
X"0177",
X"FE89",
X"FF06",
X"0177",
X"02EE",
X"02EE",
X"055F",
X"0CB2",
X"1CCF",
X"22AB",
X"101D",
X"F6B9",
X"E237",
X"DCD8",
X"E2B4",
X"EB7E",
X"F4C5",
X"FF06",
X"0B3B",
X"0F23",
X"0BB8",
X"06D6",
X"036B",
X"0000",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FD8F",
X"FC95",
X"FD12",
X"007D",
X"00FA",
X"FE89",
X"FE0C",
X"007D",
X"03E8",
X"04E2",
X"05DC",
X"0A41",
X"19E1",
X"2599",
X"1482",
X"F9A7",
X"E4A8",
X"DC5B",
X"E237",
X"EA07",
X"F254",
X"FC95",
X"0A41",
X"109A",
X"0DAC",
X"084D",
X"036B",
X"0000",
X"FD12",
X"FD12",
X"FE0C",
X"FD8F",
X"FC95",
X"FC18",
X"FD12",
X"FF83",
X"00FA",
X"FF06",
X"FE89",
X"00FA",
X"036B",
X"04E2",
X"0659",
X"0947",
X"157C",
X"249F",
X"1964",
X"FE89",
X"E98A",
X"DECC",
X"E13D",
X"E890",
X"F060",
X"F8AD",
X"0753",
X"101D",
X"0E29",
X"08CA",
X"03E8",
X"0000",
X"FC95",
X"FC18",
X"FD12",
X"FF06",
X"FD8F",
X"FC18",
X"FC18",
X"FD8F",
X"FF83",
X"FE89",
X"FE89",
X"00FA",
X"03E8",
X"0659",
X"0659",
X"084D",
X"1194",
X"222E",
X"1F40",
X"05DC",
X"EDEF",
X"DF49",
X"DF49",
X"E69C",
X"EEE9",
X"F6B9",
X"036B",
X"0EA6",
X"0EA6",
X"09C4",
X"03E8",
X"0000",
X"FD12",
X"FC95",
X"FD8F",
X"0000",
X"0000",
X"FE0C",
X"FB9B",
X"FB9B",
X"FF06",
X"FF06",
X"FE89",
X"0000",
X"0177",
X"04E2",
X"0753",
X"08CA",
X"0FA0",
X"1EC3",
X"21B1",
X"0A41",
X"F0DD",
X"E043",
X"DE4F",
X"E5A2",
X"EDEF",
X"F6B9",
X"0271",
X"0E29",
X"0E29",
X"08CA",
X"03E8",
X"007D",
X"FC95",
X"FB1E",
X"FC95",
X"FF06",
X"007D",
X"FF06",
X"FD12",
X"FC95",
X"FE89",
X"FE0C",
X"FD12",
X"FF06",
X"0271",
X"06D6",
X"08CA",
X"08CA",
X"0B3B",
X"18E7",
X"249F",
X"1388",
X"F8AD",
X"E42B",
X"DCD8",
X"E1BA",
X"EA07",
X"F2D1",
X"FE0C",
X"0CB2",
X"109A",
X"0B3B",
X"05DC",
X"0177",
X"FD8F",
X"FB9B",
X"FC95",
X"FE0C",
X"007D",
X"FF06",
X"FD8F",
X"FC95",
X"FD12",
X"FE0C",
X"FD12",
X"FE0C",
X"FF83",
X"0271",
X"0659",
X"08CA",
X"0B3B",
X"157C",
X"249F",
X"1ADB",
X"00FA",
X"E90D",
X"DCD8",
X"E0C0",
X"E98A",
X"F15A",
X"F9A7",
X"084D",
X"101D",
X"0CB2",
X"0659",
X"0271",
X"FE89",
X"FB1E",
X"FB1E",
X"FD12",
X"0000",
X"007D",
X"FE89",
X"FD8F",
X"FE0C",
X"FF83",
X"FD12",
X"FC18",
X"FE0C",
X"007D",
X"0465",
X"07D0",
X"0B3B",
X"1482",
X"23A5",
X"1D4C",
X"03E8",
X"EBFB",
X"DE4F",
X"E043",
X"E90D",
X"F15A",
X"F830",
X"055F",
X"101D",
X"0EA6",
X"084D",
X"036B",
X"FE89",
X"FAA1",
X"FAA1",
X"FD12",
X"007D",
X"0177",
X"007D",
X"FE89",
X"FE0C",
X"FE89",
X"FC18",
X"FAA1",
X"FC18",
X"FE0C",
X"0177",
X"05DC",
X"0BB8",
X"157C",
X"249F",
X"1FBD",
X"0659",
X"EDEF",
X"DF49",
X"DFC6",
X"E796",
X"F060",
X"F830",
X"0465",
X"0FA0",
X"101D",
X"09C4",
X"03E8",
X"FE89",
X"F9A7",
X"F9A7",
X"FC95",
X"FF83",
X"0177",
X"0177",
X"0000",
X"FF83",
X"FF83",
X"FC18",
X"F9A7",
X"FB1E",
X"FD8F",
X"00FA",
X"04E2",
X"0B3B",
X"1676",
X"2599",
X"1F40",
X"04E2",
X"ED72",
X"DECC",
X"E043",
X"E69C",
X"EEE9",
X"F830",
X"06D6",
X"1117",
X"109A",
X"0ABE",
X"04E2",
X"FE0C",
X"F830",
X"F736",
X"FAA1",
X"FE0C",
X"00FA",
X"01F4",
X"0177",
X"00FA",
X"FF83",
X"FB9B",
X"F9A7",
X"FB1E",
X"FD8F",
X"007D",
X"055F",
X"0CB2",
X"186A",
X"280A",
X"1FBD",
X"04E2",
X"EB7E",
X"DCD8",
X"DE4F",
X"E5A2",
X"ECF5",
X"F7B3",
X"08CA",
X"1482",
X"1388",
X"0D2F",
X"0659",
X"FE0C",
X"F736",
X"F542",
X"F7B3",
X"FC18",
X"0000",
X"0271",
X"02EE",
X"01F4",
X"0000",
X"FB9B",
X"F92A",
X"FAA1",
X"FD12",
X"007D",
X"05DC",
X"0E29",
X"1ADB",
X"2887",
X"1EC3",
X"0271",
X"EA07",
X"DC5B",
X"DECC",
X"E61F",
X"EE6C",
X"F830",
X"0947",
X"1482",
X"1388",
X"0DAC",
X"05DC",
X"FD8F",
X"F6B9",
X"F4C5",
X"F7B3",
X"FC18",
X"007D",
X"02EE",
X"02EE",
X"01F4",
X"00FA",
X"FC18",
X"F8AD",
X"F92A",
X"FB1E",
X"FF06",
X"05DC",
X"0F23",
X"1BD5",
X"2887",
X"1D4C",
X"0177",
X"EA07",
X"DD55",
X"DF49",
X"E61F",
X"EE6C",
X"F92A",
X"09C4",
X"1482",
X"128E",
X"0C35",
X"055F",
X"FE89",
X"F830",
X"F63C",
X"F7B3",
X"FD12",
X"00FA",
X"01F4",
X"0177",
X"00FA",
X"01F4",
X"FE0C",
X"F92A",
X"F830",
X"F9A7",
X"FF06",
X"06D6",
X"101D",
X"1DC9",
X"278D",
X"186A",
X"FD8F",
X"E813",
X"DF49",
X"E2B4",
X"E813",
X"EF66",
X"FAA1",
X"0ABE",
X"1405",
X"1194",
X"0B3B",
X"0465",
X"FD12",
X"F736",
X"F448",
X"F736",
X"FE0C",
X"01F4",
X"036B",
X"0271",
X"0177",
X"0177",
X"FD8F",
X"F92A",
X"F830",
X"FA24",
X"FF06",
X"06D6",
X"1194",
X"21B1",
X"2710",
X"128E",
X"F7B3",
X"E42B",
X"E043",
X"E525",
X"EA07",
X"F15A",
X"FE89",
X"0DAC",
X"1405",
X"1117",
X"0B3B",
X"03E8",
X"FC18",
X"F6B9",
X"F542",
X"F7B3",
X"FD12",
X"0000",
X"0271",
X"02EE",
X"0177",
X"007D",
X"FD8F",
X"FAA1",
X"F9A7",
X"FB1E",
X"0000",
X"07D0",
X"1405",
X"249F",
X"2328",
X"0B3B",
X"F0DD",
X"E1BA",
X"E331",
X"E890",
X"ECF5",
X"F3CB",
X"0271",
X"101D",
X"130B",
X"0FA0",
X"0947",
X"01F4",
X"FAA1",
X"F5BF",
X"F542",
X"F830",
X"FD12",
X"007D",
X"01F4",
X"01F4",
X"0177",
X"0000",
X"FE89",
X"FD12",
X"FD8F",
X"FD8F",
X"007D",
X"084D",
X"16F3",
X"249F",
X"19E1",
X"00FA",
X"EB01",
X"E2B4",
X"E719",
X"EBFB",
X"EF66",
X"F7B3",
X"07D0",
X"1117",
X"1194",
X"0E29",
X"084D",
X"0177",
X"FA24",
X"F5BF",
X"F542",
X"F830",
X"FC18",
X"FF06",
X"00FA",
X"01F4",
X"0177",
X"FF83",
X"FF06",
X"FF83",
X"007D",
X"007D",
X"0271",
X"0A41",
X"1C52",
X"222E",
X"0F23",
X"F736",
X"E5A2",
X"E3AE",
X"E98A",
X"EDEF",
X"F1D7",
X"FD8F",
X"0C35",
X"1117",
X"109A",
X"0DAC",
X"0753",
X"00FA",
X"FAA1",
X"F5BF",
X"F4C5",
X"F830",
X"FC18",
X"FE0C",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"02EE",
X"0465",
X"0753",
X"1194",
X"1F40",
X"19E1",
X"03E8",
X"EDEF",
X"E3AE",
X"E719",
X"EC78",
X"EFE3",
X"F542",
X"0271",
X"0DAC",
X"0FA0",
X"0E29",
X"0B3B",
X"05DC",
X"007D",
X"FAA1",
X"F6B9",
X"F6B9",
X"F9A7",
X"FC18",
X"FD8F",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"0000",
X"01F4",
X"03E8",
X"04E2",
X"07D0",
X"1405",
X"1FBD",
X"14FF",
X"FE0C",
X"EA07",
X"E3AE",
X"E90D",
X"EE6C",
X"F15A",
X"F8AD",
X"0659",
X"0F23",
X"0FA0",
X"0DAC",
X"09C4",
X"03E8",
X"FE89",
X"F92A",
X"F736",
X"F830",
X"FA24",
X"FC18",
X"FE0C",
X"FF06",
X"FE89",
X"FD8F",
X"FD8F",
X"0000",
X"0271",
X"0465",
X"0753",
X"0CB2",
X"1964",
X"1E46",
X"0E29",
X"F7B3",
X"E719",
X"E42B",
X"E90D",
X"EDEF",
X"F254",
X"FD12",
X"0ABE",
X"109A",
X"0FA0",
X"0CB2",
X"07D0",
X"0177",
X"FC95",
X"F7B3",
X"F736",
X"F9A7",
X"FC18",
X"FD8F",
X"FE0C",
X"FE89",
X"FE89",
X"FE0C",
X"FD12",
X"FF06",
X"0177",
X"055F",
X"09C4",
X"1211",
X"1FBD",
X"1C52",
X"06D6",
X"F060",
X"E331",
X"E4A8",
X"EA07",
X"EDEF",
X"F542",
X"03E8",
X"0F23",
X"109A",
X"0E29",
X"0ABE",
X"055F",
X"FF06",
X"F8AD",
X"F542",
X"F7B3",
X"FB9B",
X"FE0C",
X"FF06",
X"FF83",
X"FF83",
X"FE89",
X"FD8F",
X"FD8F",
X"FF83",
X"0177",
X"055F",
X"0BB8",
X"1964",
X"22AB",
X"14FF",
X"FD12",
X"E98A",
X"E2B4",
X"E69C",
X"EB01",
X"EF66",
X"F92A",
X"07D0",
X"0FA0",
X"109A",
X"0EA6",
X"0947",
X"0271",
X"FC95",
X"F736",
X"F542",
X"F7B3",
X"FB9B",
X"FE89",
X"0000",
X"00FA",
X"0000",
X"FE89",
X"FE0C",
X"FF83",
X"01F4",
X"02EE",
X"055F",
X"0D2F",
X"1DC9",
X"222E",
X"0E29",
X"F542",
X"E42B",
X"E237",
X"E813",
X"EBFB",
X"F15A",
X"FE0C",
X"0CB2",
X"1194",
X"109A",
X"0DAC",
X"0753",
X"0177",
X"FB9B",
X"F5BF",
X"F4C5",
X"F830",
X"FB9B",
X"FE0C",
X"FF06",
X"FF06",
X"FE0C",
X"FD8F",
X"FF06",
X"0177",
X"0465",
X"05DC",
X"084D",
X"1388",
X"2134",
X"1B58",
X"03E8",
X"ED72",
X"E237",
X"E4A8",
X"EA07",
X"EE6C",
X"F542",
X"036B",
X"0EA6",
X"1194",
X"0FA0",
X"0B3B",
X"04E2",
X"FF06",
X"FA24",
X"F63C",
X"F63C",
X"F8AD",
X"FC95",
X"FE0C",
X"FF06",
X"FF06",
X"FD8F",
X"FD12",
X"FE89",
X"01F4",
X"04E2",
X"0659",
X"09C4",
X"1676",
X"22AB",
X"16F3",
X"FE89",
X"E90D",
X"E1BA",
X"E796",
X"EBFB",
X"EF66",
X"F8AD",
X"06D6",
X"109A",
X"101D",
X"0D2F",
X"08CA",
X"03E8",
X"FF06",
X"F8AD",
X"F6B9",
X"F830",
X"FAA1",
X"FD8F",
X"FF06",
X"0000",
X"FE89",
X"FC18",
X"FC18",
X"FF06",
X"0271",
X"04E2",
X"0753",
X"0D2F",
X"1BD5",
X"21B1",
X"0FA0",
X"F736",
X"E525",
X"E237",
X"E813",
X"EC78",
X"F0DD",
X"FC95",
X"0B3B",
X"1194",
X"101D",
X"0CB2",
X"0753",
X"0271",
X"FD8F",
X"F830",
X"F6B9",
X"F8AD",
X"FB9B",
X"FD12",
X"FE0C",
X"FF06",
X"FE89",
X"FC95",
X"FC95",
X"FF83",
X"03E8",
X"0659",
X"0947",
X"1211",
X"2134",
X"1DC9",
X"0659",
X"EDEF",
X"E13D",
X"E42B",
X"EA07",
X"EDEF",
X"F542",
X"03E8",
X"0FA0",
X"1117",
X"0EA6",
X"09C4",
X"0465",
X"0000",
X"FAA1",
X"F6B9",
X"F830",
X"FC18",
X"FD8F",
X"FE0C",
X"FF06",
X"FF06",
X"FD8F",
X"FC18",
X"FC95",
X"0000",
X"03E8",
X"084D",
X"0DAC",
X"1BD5",
X"22AB",
X"1194",
X"F8AD",
X"E4A8",
X"E0C0",
X"E719",
X"ECF5",
X"F1D7",
X"FC95",
X"0B3B",
X"1194",
X"109A",
X"0E29",
X"0753",
X"007D",
X"FC18",
X"F6B9",
X"F5BF",
X"F92A",
X"FB9B",
X"FD8F",
X"FF83",
X"00FA",
X"FF83",
X"FD12",
X"FB9B",
X"FD12",
X"0177",
X"055F",
X"09C4",
X"1117",
X"1FBD",
X"203A",
X"0B3B",
X"F254",
X"E13D",
X"E13D",
X"E813",
X"ED72",
X"F3CB",
X"007D",
X"0EA6",
X"1211",
X"109A",
X"0D2F",
X"0659",
X"007D",
X"FAA1",
X"F63C",
X"F736",
X"FAA1",
X"FC18",
X"FD12",
X"FF83",
X"FF83",
X"FD12",
X"FAA1",
X"FAA1",
X"FF06",
X"036B",
X"0753",
X"0DAC",
X"18E7",
X"249F",
X"19E1",
X"00FA",
X"E90D",
X"DE4F",
X"E1BA",
X"E719",
X"ED72",
X"F736",
X"0753",
X"130B",
X"1482",
X"1211",
X"0CB2",
X"04E2",
X"FE0C",
X"F830",
X"F448",
X"F5BF",
X"F9A7",
X"FD12",
X"FE89",
X"FF06",
X"FE89",
X"FD12",
X"FB1E",
X"FB1E",
X"FE89",
X"036B",
X"08CA",
X"0FA0",
X"1B58",
X"249F",
X"1676",
X"FD12",
X"E796",
X"DF49",
X"E2B4",
X"E796",
X"EDEF",
X"FA24",
X"0ABE",
X"1405",
X"1388",
X"101D",
X"0947",
X"01F4",
X"FC18",
X"F736",
X"F542",
X"F830",
X"FD12",
X"FF06",
X"0000",
X"0000",
X"FD8F",
X"FA24",
X"F8AD",
X"FB1E",
X"0000",
X"04E2",
X"0BB8",
X"14FF",
X"251C",
X"251C",
X"0BB8",
X"F0DD",
X"DFC6",
X"DF49",
X"E42B",
X"E90D",
X"EF66",
X"007D",
X"1117",
X"1482",
X"130B",
X"0F23",
X"08CA",
X"0177",
X"FAA1",
X"F5BF",
X"F5BF",
X"F9A7",
X"FC18",
X"FD8F",
X"FF06",
X"FF83",
X"FD12",
X"FA24",
X"F9A7",
X"FE0C",
X"02EE",
X"0659",
X"0C35",
X"186A",
X"2616",
X"1CCF",
X"02EE",
X"EA84",
X"DE4F",
X"E13D",
X"E61F",
X"EB7E",
X"F63C",
X"084D",
X"1388",
X"1482",
X"1194",
X"0BB8",
X"0465",
X"FE0C",
X"F830",
X"F542",
X"F736",
X"FB9B",
X"FE0C",
X"FF06",
X"FF83",
X"FF06",
X"FC18",
X"FA24",
X"FA24",
X"FE89",
X"036B",
X"07D0",
X"0E29",
X"1C52",
X"2616",
X"15F9",
X"FB9B",
X"E61F",
X"DF49",
X"E331",
X"E796",
X"ECF5",
X"FA24",
X"0C35",
X"1482",
X"1405",
X"109A",
X"0ABE",
X"02EE",
X"FD12",
X"F736",
X"F5BF",
X"F8AD",
X"FB1E",
X"FD12",
X"FE89",
X"FF83",
X"FD12",
X"FAA1",
X"FA24",
X"FD12",
X"0271",
X"05DC",
X"09C4",
X"128E",
X"22AB",
X"22AB",
X"0C35",
X"F15A",
X"DF49",
X"DE4F",
X"E42B",
X"E98A",
X"F254",
X"02EE",
X"1117",
X"1482",
X"128E",
X"0EA6",
X"07D0",
X"00FA",
X"FB1E",
X"F736",
X"F6B9",
X"F92A",
X"FC18",
X"FD8F",
X"FE89",
X"FD8F",
X"FB1E",
X"FA24",
X"FC18",
X"007D",
X"03E8",
X"06D6",
X"0A41",
X"1482",
X"2422",
X"1E46",
X"0465",
X"EB7E",
X"DFC6",
X"E1BA",
X"E69C",
X"EA84",
X"F448",
X"055F",
X"1211",
X"1482",
X"128E",
X"0E29",
X"05DC",
X"FE89",
X"F9A7",
X"F736",
X"F830",
X"F9A7",
X"FC18",
X"FE89",
X"0000",
X"FE0C",
X"FB1E",
X"F92A",
X"FC18",
X"0177",
X"04E2",
X"0753",
X"09C4",
X"15F9",
X"2422",
X"1A5E",
X"007D",
X"E98A",
X"DFC6",
X"E2B4",
X"E813",
X"ED72",
X"F8AD",
X"08CA",
X"109A",
X"1194",
X"1194",
X"0D2F",
X"055F",
X"FF06",
X"FA24",
X"F830",
X"F7B3",
X"F7B3",
X"F92A",
X"FC18",
X"FE0C",
X"FE0C",
X"FC18",
X"FB1E",
X"FE89",
X"0271",
X"055F",
X"0947",
X"0DAC",
X"1B58",
X"2422",
X"1388",
X"F8AD",
X"E4A8",
X"DF49",
X"E3AE",
X"E90D",
X"EE6C",
X"FB9B",
X"0C35",
X"1388",
X"1388",
X"1117",
X"0ABE",
X"03E8",
X"FD12",
X"F736",
X"F4C5",
X"F6B9",
X"F9A7",
X"FC95",
X"FD8F",
X"FD8F",
X"FD8F",
X"FC95",
X"FD8F",
X"007D",
X"02EE",
X"04E2",
X"084D",
X"0F23",
X"1DC9",
X"21B1",
X"0D2F",
X"F448",
X"E4A8",
X"E237",
X"E5A2",
X"E90D",
X"EFE3",
X"FF83",
X"0EA6",
X"1405",
X"1388",
X"109A",
X"09C4",
X"02EE",
X"FC95",
X"F736",
X"F542",
X"F736",
X"F9A7",
X"FC18",
X"FD8F",
X"FE0C",
X"FD12",
X"FB9B",
X"FC18",
X"007D",
X"03E8",
X"05DC",
X"084D",
X"0FA0",
X"1EC3",
X"203A",
X"0ABE",
X"F1D7",
X"E237",
X"E043",
X"E5A2",
X"EA84",
X"F2D1",
X"0271",
X"0F23",
X"1405",
X"1405",
X"109A",
X"09C4",
X"0177",
X"FA24",
X"F63C",
X"F63C",
X"F8AD",
X"FAA1",
X"FC95",
X"FE0C",
X"FE0C",
X"FE0C",
X"FC18",
X"FD12",
X"00FA",
X"03E8",
X"055F",
X"084D",
X"101D",
X"1FBD",
X"1EC3",
X"084D",
X"F060",
X"E2B4",
X"E1BA",
X"E5A2",
X"E98A",
X"F254",
X"02EE",
X"109A",
X"1482",
X"1405",
X"101D",
X"08CA",
X"0177",
X"F9A7",
X"F4C5",
X"F542",
X"F830",
X"FA24",
X"FB9B",
X"FD12",
X"FE0C",
X"FD8F",
X"FD12",
X"FE89",
X"02EE",
X"055F",
X"0753",
X"0ABE",
X"1482",
X"222E",
X"1A5E",
X"00FA",
X"E98A",
X"DFC6",
X"E1BA",
X"E69C",
X"EB7E",
X"F6B9",
X"084D",
X"1405",
X"15F9",
X"1482",
X"0F23",
X"06D6",
X"FF06",
X"F7B3",
X"F3CB",
X"F4C5",
X"F7B3",
X"FA24",
X"FC18",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"0000",
X"03E8",
X"0659",
X"08CA",
X"0BB8",
X"17ED",
X"222E",
X"157C",
X"FB1E",
X"E61F",
X"DFC6",
X"E3AE",
X"E813",
X"EC78",
X"F92A",
X"0A41",
X"1482",
X"16F3",
X"14FF",
X"0E29",
X"04E2",
X"FC18",
X"F6B9",
X"F542",
X"F6B9",
X"F8AD",
X"FAA1",
X"FC18",
X"FD8F",
X"FD8F",
X"FD12",
X"FD8F",
X"007D",
X"03E8",
X"05DC",
X"084D",
X"0C35",
X"1A5E",
X"22AB",
X"130B",
X"F830",
X"E42B",
X"DF49",
X"E42B",
X"E90D",
X"EE6C",
X"FC95",
X"0CB2",
X"14FF",
X"157C",
X"1211",
X"0BB8",
X"036B",
X"FB1E",
X"F63C",
X"F542",
X"F7B3",
X"FA24",
X"FB9B",
X"FC95",
X"FD12",
X"FD12",
X"FC95",
X"FD12",
X"00FA",
X"04E2",
X"06D6",
X"084D",
X"0CB2",
X"1B58",
X"22AB",
X"1211",
X"F6B9",
X"E2B4",
X"DDD2",
X"E331",
X"E813",
X"EEE9",
X"FE0C",
X"0F23",
X"1676",
X"15F9",
X"1194",
X"0ABE",
X"0271",
X"FA24",
X"F4C5",
X"F448",
X"F736",
X"FA24",
X"FC18",
X"FD12",
X"FE0C",
X"FE0C",
X"FD12",
X"FE89",
X"02EE",
X"06D6",
X"084D",
X"09C4",
X"0D2F",
X"1A5E",
X"1E46",
X"0D2F",
X"F3CB",
X"E1BA",
X"DECC",
X"E42B",
X"E90D",
X"F0DD",
X"007D",
X"109A",
X"1770",
X"1676",
X"1194",
X"0A41",
X"00FA",
X"F830",
X"F448",
X"F4C5",
X"F736",
X"F9A7",
X"FA24",
X"FB1E",
X"FD12",
X"FD8F",
X"FD8F",
X"0000",
X"04E2",
X"084D",
X"0947",
X"0A41",
X"0FA0",
X"1CCF",
X"1D4C",
X"09C4",
X"EEE9",
X"DF49",
X"DECC",
X"E4A8",
X"EA07",
X"F3CB",
X"0465",
X"1211",
X"16F3",
X"157C",
X"1117",
X"09C4",
X"FF83",
X"F736",
X"F3CB",
X"F542",
X"F7B3",
X"F92A",
X"FA24",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"0000",
X"05DC",
X"084D",
X"0947",
X"0ABE",
X"1117",
X"1DC9",
X"1CCF",
X"084D",
X"EDEF",
X"DF49",
X"DFC6",
X"E525",
X"EB01",
X"F448",
X"055F",
X"1388",
X"186A",
X"15F9",
X"0FA0",
X"07D0",
X"FE89",
X"F736",
X"F448",
X"F5BF",
X"F830",
X"FA24",
X"FAA1",
X"FAA1",
X"FB9B",
X"FC95",
X"FD12",
X"0000",
X"0465",
X"06D6",
X"0753",
X"084D",
X"0E29",
X"1ADB",
X"1E46",
X"0CB2",
X"F34E",
X"E331",
X"E0C0",
X"E4A8",
X"E98A",
X"F2D1",
X"02EE",
X"1194",
X"16F3",
X"1482",
X"0FA0",
X"08CA",
X"FF83",
X"F7B3",
X"F542",
X"F63C",
X"F7B3",
X"FA24",
X"FB9B",
X"FC18",
X"FD12",
X"FD12",
X"FD12",
X"FF83",
X"02EE",
X"0465",
X"055F",
X"06D6",
X"0BB8",
X"16F3",
X"1FBD",
X"1482",
X"FC95",
X"E98A",
X"E13D",
X"E331",
X"E813",
X"EFE3",
X"FD8F",
X"0CB2",
X"1482",
X"130B",
X"0FA0",
X"09C4",
X"0177",
X"F92A",
X"F5BF",
X"F5BF",
X"F7B3",
X"FAA1",
X"FB9B",
X"FC95",
X"FE89",
X"FF06",
X"FE89",
X"007D",
X"0271",
X"036B",
X"02EE",
X"04E2",
X"0A41",
X"14FF",
X"1EC3",
X"157C",
X"FE89",
X"EB01",
X"E1BA",
X"E3AE",
X"E90D",
X"F060",
X"FC95",
X"0BB8",
X"1388",
X"130B",
X"0F23",
X"0947",
X"0177",
X"F9A7",
X"F63C",
X"F5BF",
X"F830",
X"FB1E",
X"FC95",
X"FC95",
X"FE0C",
X"FF83",
X"FF06",
X"0000",
X"0177",
X"01F4",
X"0271",
X"055F",
X"0BB8",
X"15F9",
X"1EC3",
X"1482",
X"FD12",
X"EA07",
X"E237",
X"E4A8",
X"EA84",
X"F1D7",
X"FE0C",
X"0CB2",
X"1388",
X"1211",
X"0E29",
X"07D0",
X"FF06",
X"F830",
X"F5BF",
X"F63C",
X"F8AD",
X"FC18",
X"FD12",
X"FD12",
X"FE0C",
X"FF83",
X"FF83",
X"0000",
X"01F4",
X"0271",
X"02EE",
X"04E2",
X"0ABE",
X"14FF",
X"1C52",
X"1388",
X"FD8F",
X"EBFB",
X"E3AE",
X"E5A2",
X"EB01",
X"F254",
X"FD8F",
X"0BB8",
X"1388",
X"128E",
X"0EA6",
X"0753",
X"FF06",
X"F830",
X"F542",
X"F5BF",
X"F830",
X"FB9B",
X"FD8F",
X"FD8F",
X"FE89",
X"007D",
X"007D",
X"007D",
X"0177",
X"01F4",
X"0177",
X"02EE",
X"0947",
X"130B",
X"1C52",
X"157C",
X"00FA",
X"EE6C",
X"E525",
X"E5A2",
X"EA07",
X"F060",
X"FB9B",
X"09C4",
X"128E",
X"128E",
X"0E29",
X"084D",
X"007D",
X"F9A7",
X"F5BF",
X"F5BF",
X"F830",
X"FB1E",
X"FC95",
X"FD12",
X"FE89",
X"00FA",
X"0177",
X"0177",
X"0271",
X"0177",
X"0000",
X"0177",
X"0753",
X"109A",
X"1964",
X"1770",
X"05DC",
X"F448",
X"E813",
X"E5A2",
X"E98A",
X"EEE9",
X"F8AD",
X"055F",
X"101D",
X"128E",
X"0F23",
X"0947",
X"01F4",
X"FAA1",
X"F6B9",
X"F63C",
X"F7B3",
X"FA24",
X"FC95",
X"FE0C",
X"FF83",
X"0177",
X"00FA",
X"0177",
X"01F4",
X"007D",
X"FF06",
X"0177",
X"07D0",
X"101D",
X"186A",
X"1676",
X"0753",
X"F5BF",
X"E90D",
X"E69C",
X"EA07",
X"EFE3",
X"F8AD",
X"0465",
X"0E29",
X"1117",
X"0DAC",
X"084D",
X"0177",
X"FB1E",
X"F736",
X"F63C",
X"F830",
X"FAA1",
X"FD12",
X"FE0C",
X"FF83",
X"00FA",
X"0177",
X"0177",
X"0177",
X"007D",
X"007D",
X"03E8",
X"0A41",
X"128E",
X"186A",
X"130B",
X"01F4",
X"F1D7",
X"E796",
X"E719",
X"EB7E",
X"F1D7",
X"FB9B",
X"06D6",
X"0F23",
X"1117",
X"0DAC",
X"07D0",
X"007D",
X"F9A7",
X"F63C",
X"F5BF",
X"F830",
X"FB9B",
X"FD8F",
X"FE89",
X"FF83",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"00FA",
X"04E2",
X"0BB8",
X"14FF",
X"19E1",
X"1117",
X"FF06",
X"EE6C",
X"E69C",
X"E813",
X"ECF5",
X"F3CB",
X"FD12",
X"084D",
X"101D",
X"109A",
X"0D2F",
X"0659",
X"FE89",
X"F92A",
X"F6B9",
X"F6B9",
X"F92A",
X"FC18",
X"FD8F",
X"FE0C",
X"FE89",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"01F4",
X"05DC",
X"0D2F",
X"15F9",
X"1964",
X"0E29",
X"FB1E",
X"EBFB",
X"E69C",
X"E90D",
X"EDEF",
X"F542",
X"FF06",
X"09C4",
X"101D",
X"101D",
X"0C35",
X"05DC",
X"FE0C",
X"F8AD",
X"F63C",
X"F736",
X"FAA1",
X"FC95",
X"FD8F",
X"FD8F",
X"FE89",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"02EE",
X"06D6",
X"0E29",
X"1770",
X"17ED",
X"09C4",
X"F736",
X"EA84",
X"E813",
X"EB7E",
X"EFE3",
X"F6B9",
X"0177",
X"0BB8",
X"101D",
X"0F23",
X"0B3B",
X"03E8",
X"FC95",
X"F736",
X"F542",
X"F736",
X"FB1E",
X"FD8F",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"036B",
X"084D",
X"1117",
X"1964",
X"157C",
X"03E8",
X"F1D7",
X"E890",
X"E90D",
X"ECF5",
X"F0DD",
X"F8AD",
X"0465",
X"0DAC",
X"109A",
X"0EA6",
X"0A41",
X"02EE",
X"FB1E",
X"F5BF",
X"F448",
X"F6B9",
X"FB9B",
X"FE0C",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"0177",
X"0271",
X"04E2",
X"0A41",
X"1388",
X"18E7",
X"109A",
X"FE89",
X"EF66",
X"E90D",
X"EA07",
X"ED72",
X"F254",
X"FB9B",
X"0753",
X"0E29",
X"101D",
X"0E29",
X"0947",
X"0177",
X"FA24",
X"F542",
X"F3CB",
X"F6B9",
X"FB1E",
X"FE0C",
X"FF83",
X"007D",
X"007D",
X"0000",
X"FF83",
X"0000",
X"00FA",
X"0271",
X"055F",
X"0CB2",
X"15F9",
X"18E7",
X"0D2F",
X"FB1E",
X"ECF5",
X"E890",
X"EB01",
X"EEE9",
X"F4C5",
X"FE89",
X"08CA",
X"0EA6",
X"0FA0",
X"0CB2",
X"06D6",
X"FF83",
X"F92A",
X"F5BF",
X"F5BF",
X"F830",
X"FB9B",
X"FE0C",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"01F4",
X"03E8",
X"08CA",
X"109A",
X"17ED",
X"1482",
X"055F",
X"F448",
X"EA07",
X"E98A",
X"ECF5",
X"F15A",
X"F8AD",
X"0271",
X"0B3B",
X"0EA6",
X"0EA6",
X"0ABE",
X"0465",
X"FD8F",
X"F830",
X"F5BF",
X"F6B9",
X"FA24",
X"FD12",
X"FF06",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF83",
X"0000",
X"01F4",
X"055F",
X"0BB8",
X"1482",
X"18E7",
X"0FA0",
X"FE0C",
X"EEE9",
X"E890",
X"EA07",
X"EE6C",
X"F448",
X"FC18",
X"05DC",
X"0C35",
X"0EA6",
X"0DAC",
X"084D",
X"01F4",
X"FC95",
X"F8AD",
X"F736",
X"F830",
X"FAA1",
X"FD12",
X"FF06",
X"FF83",
X"FE89",
X"FD8F",
X"FD8F",
X"FF06",
X"0271",
X"0659",
X"0ABE",
X"1194",
X"186A",
X"1405",
X"03E8",
X"F254",
X"E813",
X"E813",
X"EC78",
X"F1D7",
X"F8AD",
X"02EE",
X"0ABE",
X"0E29",
X"0E29",
X"0B3B",
X"055F",
X"FF83",
X"FA24",
X"F736",
X"F736",
X"F92A",
X"FB9B",
X"FD12",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF83",
X"0271",
X"0659",
X"0ABE",
X"109A",
X"1770",
X"157C",
X"0753",
X"F5BF",
X"E90D",
X"E69C",
X"EA84",
X"EFE3",
X"F6B9",
X"007D",
X"0A41",
X"0EA6",
X"0F23",
X"0CB2",
X"0753",
X"0177",
X"FC95",
X"F8AD",
X"F736",
X"F8AD",
X"FAA1",
X"FB9B",
X"FC95",
X"FD8F",
X"FD8F",
X"FD8F",
X"FF06",
X"01F4",
X"0659",
X"0ABE",
X"0F23",
X"14FF",
X"16F3",
X"0D2F",
X"FC18",
X"ED72",
X"E69C",
X"E813",
X"ECF5",
X"F3CB",
X"FC95",
X"0659",
X"0D2F",
X"0F23",
X"0E29",
X"0A41",
X"03E8",
X"FF06",
X"FB1E",
X"F8AD",
X"F8AD",
X"FA24",
X"FB9B",
X"FC18",
X"FC95",
X"FC18",
X"FB9B",
X"FC18",
X"FE89",
X"036B",
X"08CA",
X"0DAC",
X"130B",
X"18E7",
X"15F9",
X"07D0",
X"F63C",
X"E890",
X"E4A8",
X"E813",
X"EE6C",
X"F63C",
X"007D",
X"09C4",
X"0EA6",
X"0FA0",
X"0CB2",
X"0753",
X"0177",
X"FD8F",
X"FA24",
X"F8AD",
X"FA24",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FB1E",
X"FB1E",
X"FC95",
X"0000",
X"055F",
X"0ABE",
X"1117",
X"17ED",
X"1ADB",
X"1117",
X"FF06",
X"EDEF",
X"E525",
X"E5A2",
X"EA07",
X"F15A",
X"FAA1",
X"05DC",
X"0E29",
X"101D",
X"0E29",
X"09C4",
X"036B",
X"FE89",
X"FB9B",
X"F92A",
X"F92A",
X"FB1E",
X"FC95",
X"FD8F",
X"FD8F",
X"FC18",
X"FAA1",
X"FAA1",
X"FD12",
X"01F4",
X"07D0",
X"0EA6",
X"15F9",
X"1ADB",
X"15F9",
X"06D6",
X"F448",
X"E719",
X"E3AE",
X"E69C",
X"ED72",
X"F63C",
X"00FA",
X"0B3B",
X"101D",
X"109A",
X"0DAC",
X"0753",
X"01F4",
X"FD8F",
X"FAA1",
X"F92A",
X"FA24",
X"FB9B",
X"FC95",
X"FC95",
X"FC18",
X"FB1E",
X"FA24",
X"FAA1",
X"FE0C",
X"04E2",
X"0C35",
X"1388",
X"1A5E",
X"1B58",
X"0FA0",
X"FD12",
X"EB01",
X"E2B4",
X"E4A8",
X"EA07",
X"F15A",
X"FB1E",
X"06D6",
X"0F23",
X"1194",
X"0FA0",
X"0ABE",
X"055F",
X"0000",
X"FC18",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FB9B",
X"FB1E",
X"FA24",
X"FAA1",
X"FC95",
X"0177",
X"07D0",
X"0FA0",
X"17ED",
X"1DC9",
X"17ED",
X"0659",
X"F1D7",
X"E42B",
X"E237",
X"E719",
X"EDEF",
X"F5BF",
X"00FA",
X"0C35",
X"1194",
X"1194",
X"0DAC",
X"0753",
X"01F4",
X"FD8F",
X"FA24",
X"F92A",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FB9B",
X"FB1E",
X"FB1E",
X"FC18",
X"FF83",
X"0465",
X"0A41",
X"1117",
X"186A",
X"1B58",
X"128E",
X"0000",
X"ED72",
X"E331",
X"E3AE",
X"E90D",
X"EFE3",
X"F8AD",
X"0465",
X"0DAC",
X"1194",
X"109A",
X"0C35",
X"06D6",
X"01F4",
X"FD12",
X"F9A7",
X"F92A",
X"FAA1",
X"FB9B",
X"FC18",
X"FC18",
X"FB1E",
X"F9A7",
X"F92A",
X"FAA1",
X"FF83",
X"05DC",
X"0D2F",
X"1482",
X"1B58",
X"1B58",
X"0F23",
X"FB1E",
X"E98A",
X"E237",
X"E42B",
X"EA07",
X"F1D7",
X"FC18",
X"07D0",
X"0FA0",
X"1117",
X"0F23",
X"09C4",
X"04E2",
X"0000",
X"FC18",
X"F9A7",
X"FA24",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FAA1",
X"F92A",
X"F92A",
X"FC18",
X"00FA",
X"0753",
X"0DAC",
X"14FF",
X"1B58",
X"19E1",
X"0C35",
X"F7B3",
X"E796",
X"E2B4",
X"E61F",
X"EC78",
X"F448",
X"FF06",
X"09C4",
X"101D",
X"109A",
X"0CB2",
X"06D6",
X"01F4",
X"FD8F",
X"FAA1",
X"FA24",
X"FB1E",
X"FD12",
X"FD8F",
X"FD12",
X"FC18",
X"FA24",
X"F8AD",
X"F92A",
X"FC95",
X"01F4",
X"084D",
X"101D",
X"17ED",
X"1CCF",
X"186A",
X"0753",
X"F1D7",
X"E3AE",
X"E1BA",
X"E796",
X"EEE9",
X"F6B9",
X"00FA",
X"0BB8",
X"1117",
X"109A",
X"0BB8",
X"0659",
X"0177",
X"FD12",
X"FAA1",
X"FA24",
X"FB9B",
X"FD12",
X"FD12",
X"FC95",
X"FB9B",
X"FA24",
X"F8AD",
X"FA24",
X"FE89",
X"0465",
X"0ABE",
X"1211",
X"1964",
X"1CCF",
X"1405",
X"007D",
X"EC78",
X"E237",
X"E2B4",
X"E890",
X"EFE3",
X"F92A",
X"0465",
X"0DAC",
X"1194",
X"101D",
X"0BB8",
X"05DC",
X"0000",
X"FC18",
X"FA24",
X"FAA1",
X"FC18",
X"FD12",
X"FD8F",
X"FC95",
X"FB1E",
X"F92A",
X"F8AD",
X"FAA1",
X"FF83",
X"0659",
X"0D2F",
X"14FF",
X"1C52",
X"1BD5",
X"0F23",
X"FA24",
X"E890",
X"E13D",
X"E3AE",
X"E98A",
X"F1D7",
X"FC18",
X"0753",
X"0FA0",
X"1211",
X"101D",
X"0ABE",
X"0465",
X"FF06",
X"FB1E",
X"FA24",
X"FAA1",
X"FC18",
X"FC95",
X"FC95",
X"FC18",
X"FB1E",
X"F9A7",
X"F92A",
X"FB9B",
X"007D",
X"06D6",
X"0DAC",
X"157C",
X"1B58",
X"1964",
X"0C35",
X"F830",
X"E90D",
X"E331",
X"E61F",
X"EBFB",
X"F3CB",
X"FE0C",
X"084D",
X"0F23",
X"101D",
X"0D2F",
X"07D0",
X"0271",
X"FE0C",
X"FB1E",
X"FAA1",
X"FC18",
X"FD8F",
X"FE0C",
X"FD8F",
X"FC18",
X"FA24",
X"F7B3",
X"F7B3",
X"FB9B",
X"01F4",
X"08CA",
X"101D",
X"17ED",
X"1D4C",
X"18E7",
X"084D",
X"F2D1",
X"E4A8",
X"E1BA",
X"E719",
X"EE6C",
X"F6B9",
X"00FA",
X"0B3B",
X"109A",
X"101D",
X"0BB8",
X"05DC",
X"00FA",
X"FC95",
X"FAA1",
X"FAA1",
X"FC18",
X"FE0C",
X"FE89",
X"FE0C",
X"FC18",
X"F92A",
X"F736",
X"F830",
X"FC95",
X"02EE",
X"0A41",
X"1211",
X"19E1",
X"1D4C",
X"157C",
X"02EE",
X"EE6C",
X"E2B4",
X"E1BA",
X"E813",
X"F060",
X"FA24",
X"04E2",
X"0DAC",
X"1117",
X"0FA0",
X"0ABE",
X"0465",
X"FF06",
X"FAA1",
X"F9A7",
X"FB1E",
X"FD12",
X"FE89",
X"FF06",
X"FD8F",
X"FB9B",
X"F8AD",
X"F7B3",
X"F92A",
X"FD8F",
X"0465",
X"0B3B",
X"1405",
X"1CCF",
X"1E46",
X"1211",
X"FD12",
X"EA07",
X"E13D",
X"E331",
X"E90D",
X"F15A",
X"FC18",
X"084D",
X"101D",
X"128E",
X"0FA0",
X"0947",
X"02EE",
X"FD12",
X"F92A",
X"F8AD",
X"FA24",
X"FD12",
X"FF06",
X"FF06",
X"FD8F",
X"FB1E",
X"F92A",
X"F92A",
X"FB1E",
X"FF06",
X"055F",
X"0CB2",
X"157C",
X"1D4C",
X"1CCF",
X"0E29",
X"F92A",
X"E813",
X"E237",
X"E42B",
X"EA07",
X"F2D1",
X"FE89",
X"09C4",
X"101D",
X"109A",
X"0CB2",
X"06D6",
X"00FA",
X"FC95",
X"FAA1",
X"FAA1",
X"FC18",
X"FE89",
X"FF83",
X"FE89",
X"FC95",
X"FA24",
X"F830",
X"F9A7",
X"FD8F",
X"01F4",
X"0753",
X"0D2F",
X"14FF",
X"1CCF",
X"1A5E",
X"09C4",
X"F4C5",
X"E5A2",
X"E237",
X"E5A2",
X"EBFB",
X"F542",
X"0177",
X"0CB2",
X"1194",
X"1117",
X"0CB2",
X"0659",
X"0000",
X"FB9B",
X"F92A",
X"F92A",
X"FB1E",
X"FD12",
X"FE0C",
X"FE0C",
X"FC95",
X"FB1E",
X"FA24",
X"FC18",
X"FF83",
X"03E8",
X"07D0",
X"0CB2",
X"1388",
X"1B58",
X"186A",
X"08CA",
X"F448",
X"E69C",
X"E331",
X"E69C",
X"ECF5",
X"F5BF",
X"01F4",
X"0BB8",
X"101D",
X"0FA0",
X"0C35",
X"0659",
X"00FA",
X"FC95",
X"F9A7",
X"F92A",
X"FB1E",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FB1E",
X"FB1E",
X"FC95",
X"FF83",
X"02EE",
X"0753",
X"0D2F",
X"1482",
X"1C52",
X"186A",
X"0753",
X"F34E",
X"E525",
X"E2B4",
X"E719",
X"ECF5",
X"F5BF",
X"01F4",
X"0CB2",
X"1194",
X"109A",
X"0C35",
X"055F",
X"FF83",
X"FB1E",
X"F830",
X"F7B3",
X"FA24",
X"FD12",
X"FE0C",
X"FD8F",
X"FC95",
X"FC18",
X"FC18",
X"FE0C",
X"007D",
X"03E8",
X"0753",
X"0BB8",
X"1211",
X"19E1",
X"16F3",
X"0659",
X"F2D1",
X"E61F",
X"E42B",
X"E796",
X"ED72",
X"F6B9",
X"036B",
X"0DAC",
X"1117",
X"0F23",
X"0ABE",
X"0465",
X"FE89",
X"FB1E",
X"F8AD",
X"F92A",
X"FB9B",
X"FD8F",
X"FE0C",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FF06",
X"01F4",
X"0465",
X"0753",
X"0B3B",
X"1211",
X"19E1",
X"16F3",
X"06D6",
X"F3CB",
X"E61F",
X"E3AE",
X"E69C",
X"ECF5",
X"F736",
X"04E2",
X"0F23",
X"1211",
X"101D",
X"0BB8",
X"055F",
X"FE89",
X"FA24",
X"F7B3",
X"F830",
X"FA24",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FD12",
X"FD8F",
X"0000",
X"02EE",
X"05DC",
X"084D",
X"0C35",
X"128E",
X"19E1",
X"15F9",
X"055F",
X"F254",
X"E5A2",
X"E2B4",
X"E69C",
X"ECF5",
X"F736",
X"0465",
X"0EA6",
X"1211",
X"1194",
X"0D2F",
X"0659",
X"FF06",
X"FA24",
X"F7B3",
X"F7B3",
X"F8AD",
X"FAA1",
X"FB9B",
X"FC18",
X"FC95",
X"FC95",
X"FE0C",
X"007D",
X"036B",
X"05DC",
X"084D",
X"0C35",
X"1194",
X"18E7",
X"17ED",
X"07D0",
X"F448",
X"E69C",
X"E331",
X"E69C",
X"EC78",
X"F5BF",
X"0271",
X"0D2F",
X"1117",
X"0FA0",
X"0BB8",
X"05DC",
X"FF83",
X"FB9B",
X"F8AD",
X"F830",
X"F92A",
X"FA24",
X"FAA1",
X"FB1E",
X"FC95",
X"FD8F",
X"FE89",
X"00FA",
X"02EE",
X"04E2",
X"0753",
X"0B3B",
X"0FA0",
X"15F9",
X"16F3",
X"0B3B",
X"F92A",
X"EA84",
X"E42B",
X"E61F",
X"EB01",
X"F3CB",
X"0000",
X"0BB8",
X"109A",
X"0FA0",
X"0C35",
X"05DC",
X"FF06",
X"FA24",
X"F830",
X"F830",
X"F9A7",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FE89",
X"FF06",
X"00FA",
X"0271",
X"02EE",
X"0465",
X"0753",
X"0CB2",
X"1388",
X"1770",
X"101D",
X"0000",
X"EFE3",
X"E69C",
X"E61F",
X"EA84",
X"F254",
X"FD12",
X"08CA",
X"0FA0",
X"101D",
X"0D2F",
X"07D0",
X"00FA",
X"FB1E",
X"F8AD",
X"F7B3",
X"F8AD",
X"FA24",
X"FB1E",
X"FC18",
X"FE0C",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"01F4",
X"0465",
X"07D0",
X"0D2F",
X"1388",
X"1770",
X"1194",
X"01F4",
X"F1D7",
X"E796",
X"E69C",
X"EB01",
X"F254",
X"FC18",
X"0753",
X"0EA6",
X"101D",
X"0CB2",
X"06D6",
X"FF83",
X"FA24",
X"F7B3",
X"F7B3",
X"F92A",
X"FB1E",
X"FD12",
X"FE0C",
X"FF06",
X"FF06",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"0271",
X"0659",
X"0C35",
X"130B",
X"16F3",
X"1194",
X"02EE",
X"F34E",
X"E90D",
X"E719",
X"EA84",
X"F15A",
X"FAA1",
X"05DC",
X"0D2F",
X"0FA0",
X"0D2F",
X"07D0",
X"0177",
X"FB9B",
X"F8AD",
X"F736",
X"F830",
X"FA24",
X"FB9B",
X"FD12",
X"FE89",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"02EE",
X"05DC",
X"0B3B",
X"1117",
X"15F9",
X"1194",
X"03E8",
X"F448",
X"E98A",
X"E796",
X"EB7E",
X"F254",
X"FC18",
X"06D6",
X"0DAC",
X"0EA6",
X"0BB8",
X"0659",
X"0000",
X"FB1E",
X"F8AD",
X"F830",
X"F9A7",
X"FB1E",
X"FC95",
X"FD12",
X"FE0C",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"00FA",
X"02EE",
X"055F",
X"09C4",
X"0FA0",
X"157C",
X"1405",
X"084D",
X"F830",
X"EB7E",
X"E69C",
X"E98A",
X"F060",
X"F9A7",
X"04E2",
X"0CB2",
X"0F23",
X"0D2F",
X"084D",
X"0177",
X"FB1E",
X"F830",
X"F7B3",
X"F8AD",
X"FB1E",
X"FC95",
X"FD8F",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"00FA",
X"036B",
X"084D",
X"0EA6",
X"14FF",
X"157C",
X"0BB8",
X"FC18",
X"EE6C",
X"E719",
X"E890",
X"EE6C",
X"F736",
X"0177",
X"0ABE",
X"0F23",
X"0EA6",
X"0A41",
X"03E8",
X"FD12",
X"F8AD",
X"F736",
X"F7B3",
X"F9A7",
X"FB9B",
X"FD8F",
X"FF06",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"007D",
X"02EE",
X"07D0",
X"0E29",
X"14FF",
X"16F3",
X"0E29",
X"FD8F",
X"EE6C",
X"E69C",
X"E796",
X"ECF5",
X"F5BF",
X"0000",
X"0A41",
X"0F23",
X"0EA6",
X"0ABE",
X"0465",
X"FD8F",
X"F92A",
X"F736",
X"F7B3",
X"FA24",
X"FB9B",
X"FD12",
X"FE0C",
X"FF83",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0271",
X"06D6",
X"0DAC",
X"1405",
X"1676",
X"0E29",
X"FF06",
X"EFE3",
X"E796",
X"E719",
X"EC78",
X"F4C5",
X"FF83",
X"09C4",
X"0F23",
X"0FA0",
X"0BB8",
X"055F",
X"FE0C",
X"F92A",
X"F736",
X"F7B3",
X"F9A7",
X"FC18",
X"FD8F",
X"FE89",
X"FF83",
X"007D",
X"0000",
X"0000",
X"0000",
X"007D",
X"02EE",
X"0753",
X"0CB2",
X"128E",
X"14FF",
X"0EA6",
X"00FA",
X"F2D1",
X"E98A",
X"E890",
X"ECF5",
X"F448",
X"FE0C",
X"07D0",
X"0DAC",
X"0E29",
X"0ABE",
X"04E2",
X"FF06",
X"FA24",
X"F7B3",
X"F7B3",
X"F92A",
X"FB1E",
X"FC95",
X"FE0C",
X"FF83",
X"007D",
X"007D",
X"00FA",
X"007D",
X"00FA",
X"02EE",
X"06D6",
X"0C35",
X"1194",
X"1388",
X"0F23",
X"02EE",
X"F5BF",
X"EBFB",
X"E90D",
X"EBFB",
X"F2D1",
X"FC18",
X"0659",
X"0CB2",
X"0DAC",
X"0B3B",
X"0659",
X"FF83",
X"FA24",
X"F736",
X"F736",
X"F92A",
X"FB1E",
X"FD12",
X"FE89",
X"0000",
X"0177",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0271",
X"0659",
X"0C35",
X"1194",
X"1405",
X"0EA6",
X"01F4",
X"F4C5",
X"EBFB",
X"E98A",
X"EC78",
X"F34E",
X"FC95",
X"0659",
X"0CB2",
X"0DAC",
X"0B3B",
X"05DC",
X"FF83",
X"F9A7",
X"F736",
X"F736",
X"F8AD",
X"FB1E",
X"FD12",
X"FE89",
X"0000",
X"00FA",
X"0177",
X"00FA",
X"007D",
X"00FA",
X"036B",
X"07D0",
X"0DAC",
X"128E",
X"130B",
X"0BB8",
X"FE89",
X"F254",
X"EB01",
X"E98A",
X"ED72",
X"F542",
X"FF06",
X"084D",
X"0DAC",
X"0EA6",
X"0BB8",
X"05DC",
X"FF06",
X"F92A",
X"F63C",
X"F63C",
X"F830",
X"FB1E",
X"FD8F",
X"FF06",
X"007D",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"0177",
X"036B",
X"084D",
X"0E29",
X"1388",
X"1211",
X"08CA",
X"FB1E",
X"EFE3",
X"EA84",
X"EB01",
X"EF66",
X"F736",
X"00FA",
X"0947",
X"0E29",
X"0E29",
X"0ABE",
X"04E2",
X"FE0C",
X"F8AD",
X"F63C",
X"F63C",
X"F8AD",
X"FB1E",
X"FD8F",
X"FF83",
X"007D",
X"0177",
X"01F4",
X"01F4",
X"0177",
X"01F4",
X"0465",
X"0947",
X"0F23",
X"130B",
X"0FA0",
X"0465",
X"F6B9",
X"EDEF",
X"EB01",
X"EC78",
X"F1D7",
X"F9A7",
X"02EE",
X"0ABE",
X"0EA6",
X"0E29",
X"0A41",
X"036B",
X"FC95",
X"F830",
X"F63C",
X"F6B9",
X"F8AD",
X"FB9B",
X"FE0C",
X"0000",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0271",
X"055F",
X"0A41",
X"101D",
X"128E",
X"0D2F",
X"00FA",
X"F448",
X"EC78",
X"EB01",
X"EDEF",
X"F3CB",
X"FB9B",
X"04E2",
X"0BB8",
X"0EA6",
X"0D2F",
X"08CA",
X"01F4",
X"FC18",
X"F830",
X"F6B9",
X"F736",
X"F9A7",
X"FC18",
X"FE89",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"01F4",
X"036B",
X"06D6",
X"0C35",
X"1117",
X"1211",
X"0ABE",
X"FE0C",
X"F1D7",
X"EB7E",
X"EB01",
X"EEE9",
X"F542",
X"FD8F",
X"05DC",
X"0C35",
X"0EA6",
X"0D2F",
X"07D0",
X"00FA",
X"FB1E",
X"F736",
X"F63C",
X"F736",
X"F9A7",
X"FC95",
X"FF06",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"02EE",
X"055F",
X"0947",
X"0EA6",
X"128E",
X"101D",
X"055F",
X"F830",
X"EDEF",
X"EA07",
X"EBFB",
X"F15A",
X"F8AD",
X"0177",
X"0947",
X"0DAC",
X"0E29",
X"0B3B",
X"055F",
X"FF06",
X"FAA1",
X"F736",
X"F63C",
X"F7B3",
X"FA24",
X"FD12",
X"FF83",
X"007D",
X"00FA",
X"00FA",
X"01F4",
X"02EE",
X"0465",
X"0753",
X"0BB8",
X"109A",
X"1194",
X"0A41",
X"FD12",
X"F15A",
X"EB01",
X"EB7E",
X"EF66",
X"F542",
X"FD8F",
X"05DC",
X"0BB8",
X"0E29",
X"0CB2",
X"084D",
X"0271",
X"FD8F",
X"F9A7",
X"F7B3",
X"F736",
X"F8AD",
X"FB1E",
X"FD12",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"02EE",
X"055F",
X"07D0",
X"0BB8",
X"101D",
X"1211",
X"0C35",
X"0000",
X"F34E",
X"EB7E",
X"EA84",
X"EDEF",
X"F34E",
X"FAA1",
X"036B",
X"0A41",
X"0D2F",
X"0D2F",
X"0A41",
X"055F",
X"007D",
X"FC18",
X"F92A",
X"F7B3",
X"F830",
X"F9A7",
X"FB1E",
X"FC95",
X"FD8F",
X"FE89",
X"007D",
X"02EE",
X"05DC",
X"0947",
X"0CB2",
X"101D",
X"1194",
X"0DAC",
X"02EE",
X"F6B9",
X"EDEF",
X"EA84",
X"EB7E",
X"F060",
X"F7B3",
X"007D",
X"07D0",
X"0C35",
X"0D2F",
X"0BB8",
X"07D0",
X"02EE",
X"FE89",
X"FB1E",
X"F92A",
X"F8AD",
X"F92A",
X"FA24",
X"FB1E",
X"FC18",
X"FD12",
X"FF06",
X"0177",
X"055F",
X"08CA",
X"0CB2",
X"101D",
X"1211",
X"0F23",
X"0659",
X"FAA1",
X"F060",
X"EB7E",
X"EB01",
X"EDEF",
X"F448",
X"FC95",
X"055F",
X"0ABE",
X"0D2F",
X"0CB2",
X"09C4",
X"055F",
X"007D",
X"FC95",
X"FA24",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FB1E",
X"FC18",
X"FD8F",
X"FF06",
X"01F4",
X"0659",
X"0ABE",
X"0EA6",
X"1211",
X"1211",
X"0C35",
X"00FA",
X"F542",
X"ECF5",
X"EA07",
X"EB7E",
X"F0DD",
X"F92A",
X"01F4",
X"0947",
X"0CB2",
X"0D2F",
X"0ABE",
X"06D6",
X"01F4",
X"FE89",
X"FB9B",
X"FA24",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC95",
X"FD8F",
X"0000",
X"03E8",
X"08CA",
X"0D2F",
X"1194",
X"1388",
X"0FA0",
X"055F",
X"F8AD",
X"EEE9",
X"EA07",
X"EA07",
X"EE6C",
X"F5BF",
X"FF06",
X"0753",
X"0BB8",
X"0DAC",
X"0CB2",
X"08CA",
X"03E8",
X"FF06",
X"FB9B",
X"F9A7",
X"F92A",
X"FA24",
X"FB1E",
X"FB9B",
X"FC18",
X"FC18",
X"FD12",
X"FF06",
X"01F4",
X"0659",
X"0ABE",
X"101D",
X"1482",
X"130B",
X"0A41",
X"FD12",
X"F15A",
X"EA84",
X"E90D",
X"EB7E",
X"F254",
X"FB1E",
X"0465",
X"0A41",
X"0DAC",
X"0DAC",
X"0ABE",
X"05DC",
X"00FA",
X"FD8F",
X"FAA1",
X"F9A7",
X"FA24",
X"FB1E",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FD12",
X"FF83",
X"036B",
X"084D",
X"0E29",
X"1405",
X"15F9",
X"0FA0",
X"036B",
X"F5BF",
X"EBFB",
X"E813",
X"E98A",
X"EEE9",
X"F7B3",
X"00FA",
X"084D",
X"0CB2",
X"0E29",
X"0C35",
X"084D",
X"036B",
X"FF06",
X"FB9B",
X"FA24",
X"FA24",
X"FB1E",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FD8F",
X"00FA",
X"05DC",
X"0BB8",
X"1211",
X"1676",
X"1388",
X"0947",
X"FB1E",
X"EF66",
X"E90D",
X"E890",
X"EBFB",
X"F3CB",
X"FD12",
X"05DC",
X"0BB8",
X"0E29",
X"0DAC",
X"0A41",
X"055F",
X"00FA",
X"FD12",
X"FB1E",
X"FAA1",
X"FAA1",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC95",
X"FF06",
X"02EE",
X"084D",
X"0E29",
X"1482",
X"15F9",
X"0FA0",
X"0271",
X"F4C5",
X"EB01",
X"E813",
X"EA07",
X"EF66",
X"F830",
X"0177",
X"0947",
X"0D2F",
X"0E29",
X"0C35",
X"07D0",
X"02EE",
X"FF06",
X"FC18",
X"FAA1",
X"FAA1",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FD12",
X"FF83",
X"0465",
X"09C4",
X"109A",
X"15F9",
X"1482",
X"0B3B",
X"FC95",
X"F060",
X"EA07",
X"E90D",
X"EC78",
X"F2D1",
X"FB9B",
X"0465",
X"0B3B",
X"0E29",
X"0DAC",
X"0A41",
X"055F",
X"00FA",
X"FD8F",
X"FB1E",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC95",
X"FC95",
X"FC18",
X"FB9B",
X"FC18",
X"FD8F",
X"00FA",
X"05DC",
X"0C35",
X"128E",
X"15F9",
X"1211",
X"06D6",
X"F8AD",
X"EDEF",
X"E90D",
X"E98A",
X"EDEF",
X"F5BF",
X"FF06",
X"0753",
X"0C35",
X"0E29",
X"0CB2",
X"084D",
X"036B",
X"FE89",
X"FB9B",
X"FAA1",
X"FAA1",
X"FB9B",
X"FC95",
X"FD8F",
X"FD12",
X"FC95",
X"FB9B",
X"FC18",
X"FE0C",
X"01F4",
X"0753",
X"0DAC",
X"1405",
X"15F9",
X"0FA0",
X"036B",
X"F542",
X"EBFB",
X"E90D",
X"EB01",
X"F060",
X"F8AD",
X"01F4",
X"0947",
X"0CB2",
X"0D2F",
X"0ABE",
X"0659",
X"00FA",
X"FD12",
X"FB1E",
X"FB1E",
X"FC18",
X"FD12",
X"FD8F",
X"FD8F",
X"FD12",
X"FB9B",
X"FAA1",
X"FB9B",
X"FE89",
X"036B",
X"09C4",
X"101D",
X"157C",
X"14FF",
X"0C35",
X"FE89",
X"F1D7",
X"EA84",
X"E98A",
X"EC78",
X"F2D1",
X"FB9B",
X"0465",
X"0A41",
X"0CB2",
X"0CB2",
X"0947",
X"0465",
X"0000",
X"FC95",
X"FB1E",
X"FB9B",
X"FC95",
X"FD8F",
X"FE89",
X"FE0C",
X"FC95",
X"FB1E",
X"FAA1",
X"FC95",
X"0000",
X"055F",
X"0B3B",
X"1194",
X"15F9",
X"130B",
X"084D",
X"FB1E",
X"EFE3",
X"EA07",
X"E98A",
X"ED72",
X"F4C5",
X"FE0C",
X"0659",
X"0B3B",
X"0D2F",
X"0C35",
X"084D",
X"02EE",
X"FE89",
X"FB9B",
X"FAA1",
X"FB1E",
X"FC95",
X"FD8F",
X"FE0C",
X"FD12",
X"FC18",
X"FB1E",
X"FB9B",
X"FE0C",
X"01F4",
X"06D6",
X"0CB2",
X"1211",
X"14FF",
X"1117",
X"0659",
X"F9A7",
X"EF66",
X"EA84",
X"EA07",
X"EE6C",
X"F5BF",
X"FF06",
X"06D6",
X"0BB8",
X"0D2F",
X"0B3B",
X"0753",
X"0271",
X"FE0C",
X"FB9B",
X"FB1E",
X"FB9B",
X"FC95",
X"FD8F",
X"FD8F",
X"FD12",
X"FB9B",
X"FB1E",
X"FC18",
X"FF06",
X"02EE",
X"07D0",
X"0D2F",
X"1211",
X"1405",
X"101D",
X"05DC",
X"F9A7",
X"EF66",
X"EA07",
X"EA07",
X"EE6C",
X"F63C",
X"0000",
X"0753",
X"0BB8",
X"0CB2",
X"0ABE",
X"06D6",
X"01F4",
X"FD8F",
X"FB1E",
X"FAA1",
X"FB1E",
X"FC95",
X"FD8F",
X"FD8F",
X"FC95",
X"FB9B",
X"FB9B",
X"FD12",
X"0000",
X"03E8",
X"084D",
X"0DAC",
X"1211",
X"1405",
X"0FA0",
X"055F",
X"F8AD",
X"EE6C",
X"E98A",
X"EA07",
X"EEE9",
X"F736",
X"007D",
X"07D0",
X"0C35",
X"0D2F",
X"0ABE",
X"0659",
X"0177",
X"FD12",
X"FB1E",
X"FA24",
X"FB1E",
X"FC18",
X"FD12",
X"FC95",
X"FC18",
X"FB1E",
X"FB9B",
X"FD8F",
X"007D",
X"0465",
X"0947",
X"0E29",
X"128E",
X"1405",
X"0F23",
X"0465",
X"F7B3",
X"ED72",
X"E98A",
X"EA84",
X"EFE3",
X"F7B3",
X"007D",
X"084D",
X"0C35",
X"0CB2",
X"0A41",
X"05DC",
X"00FA",
X"FD12",
X"FB1E",
X"FAA1",
X"FB9B",
X"FC95",
X"FD12",
X"FC95",
X"FB9B",
X"FB1E",
X"FB9B",
X"FD8F",
X"007D",
X"0465",
X"0947",
X"0E29",
X"1211",
X"1388",
X"0EA6",
X"0465",
X"F830",
X"EE6C",
X"EA07",
X"EB7E",
X"F060",
X"F830",
X"00FA",
X"084D",
X"0C35",
X"0C35",
X"09C4",
X"055F",
X"007D",
X"FD12",
X"FB1E",
X"FAA1",
X"FB9B",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FB9B",
X"FC95",
X"FE89",
X"00FA",
X"0465",
X"08CA",
X"0D2F",
X"109A",
X"1211",
X"0E29",
X"04E2",
X"F8AD",
X"EEE9",
X"EA84",
X"EB7E",
X"F060",
X"F8AD",
X"0177",
X"08CA",
X"0C35",
X"0C35",
X"0947",
X"04E2",
X"0000",
X"FC18",
X"FAA1",
X"FAA1",
X"FB9B",
X"FC95",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FF06",
X"0177",
X"0465",
X"084D",
X"0C35",
X"0FA0",
X"109A",
X"0D2F",
X"04E2",
X"FA24",
X"F060",
X"EB7E",
X"EBFB",
X"F060",
X"F830",
X"00FA",
X"084D",
X"0C35",
X"0C35",
X"09C4",
X"04E2",
X"0000",
X"FC18",
X"FA24",
X"F9A7",
X"FAA1",
X"FB9B",
X"FC95",
X"FD12",
X"FD8F",
X"FD8F",
X"FE89",
X"FF83",
X"0177",
X"03E8",
X"06D6",
X"0ABE",
X"0EA6",
X"101D",
X"0E29",
X"0659",
X"FC18",
X"F2D1",
X"ECF5",
X"EBFB",
X"EFE3",
X"F736",
X"0000",
X"0753",
X"0BB8",
X"0C35",
X"09C4",
X"055F",
X"0000",
X"FC18",
X"F9A7",
X"F9A7",
X"FAA1",
X"FB9B",
X"FC95",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FF83",
X"00FA",
X"02EE",
X"0659",
X"09C4",
X"0DAC",
X"0FA0",
X"0E29",
X"07D0",
X"FE89",
X"F542",
X"EE6C",
X"EC78",
X"EF66",
X"F63C",
X"FE89",
X"05DC",
X"0ABE",
X"0BB8",
X"09C4",
X"05DC",
X"00FA",
X"FC95",
X"FA24",
X"F9A7",
X"FAA1",
X"FB9B",
X"FD12",
X"FE0C",
X"FE89",
X"FE0C",
X"FE0C",
X"FE89",
X"FF83",
X"0177",
X"0465",
X"084D",
X"0CB2",
X"0FA0",
X"0FA0",
X"0ABE",
X"00FA",
X"F6B9",
X"EEE9",
X"EBFB",
X"EDEF",
X"F448",
X"FC95",
X"04E2",
X"0A41",
X"0C35",
X"0ABE",
X"06D6",
X"01F4",
X"FD8F",
X"FAA1",
X"FA24",
X"FAA1",
X"FB9B",
X"FD12",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FE0C",
X"FF06",
X"00FA",
X"03E8",
X"084D",
X"0CB2",
X"101D",
X"109A",
X"0BB8",
X"01F4",
X"F6B9",
X"EE6C",
X"EB7E",
X"ED72",
X"F34E",
X"FB9B",
X"03E8",
X"09C4",
X"0C35",
X"0B3B",
X"07D0",
X"02EE",
X"FE0C",
X"FB1E",
X"FA24",
X"FAA1",
X"FC18",
X"FD8F",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FD12",
X"FE89",
X"00FA",
X"0465",
X"08CA",
X"0DAC",
X"1117",
X"1194",
X"0C35",
X"01F4",
X"F63C",
X"EDEF",
X"EA84",
X"EC78",
X"F254",
X"FAA1",
X"036B",
X"0A41",
X"0CB2",
X"0C35",
X"084D",
X"036B",
X"FE89",
X"FB9B",
X"FAA1",
X"FB1E",
X"FC18",
X"FD12",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FF06",
X"0177",
X"04E2",
X"0947",
X"0DAC",
X"109A",
X"1117",
X"0C35",
X"0271",
X"F736",
X"EE6C",
X"EA84",
X"EC78",
X"F254",
X"FA24",
X"02EE",
X"0947",
X"0C35",
X"0BB8",
X"084D",
X"036B",
X"FF06",
X"FC18",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FE0C",
X"FF83",
X"0177",
X"03E8",
X"0753",
X"0BB8",
X"0F23",
X"101D",
X"0CB2",
X"03E8",
X"F9A7",
X"F0DD",
X"ECF5",
X"ED72",
X"F254",
X"F9A7",
X"01F4",
X"084D",
X"0B3B",
X"0B3B",
X"084D",
X"036B",
X"FF06",
X"FB9B",
X"FA24",
X"FAA1",
X"FB1E",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"02EE",
X"05DC",
X"09C4",
X"0D2F",
X"0F23",
X"0CB2",
X"055F",
X"FC18",
X"F3CB",
X"EEE9",
X"EE6C",
X"F254",
X"F92A",
X"00FA",
X"06D6",
X"0A41",
X"0A41",
X"07D0",
X"036B",
X"FF06",
X"FB9B",
X"FA24",
X"FA24",
X"FB1E",
X"FC18",
X"FD12",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"01F4",
X"0465",
X"084D",
X"0BB8",
X"0E29",
X"0CB2",
X"06D6",
X"FE89",
X"F63C",
X"F0DD",
X"EF66",
X"F1D7",
X"F7B3",
X"FF83",
X"05DC",
X"09C4",
X"0A41",
X"07D0",
X"03E8",
X"FF83",
X"FC18",
X"FA24",
X"F9A7",
X"FAA1",
X"FC18",
X"FD12",
X"FE89",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"0177",
X"036B",
X"0659",
X"0A41",
X"0CB2",
X"0C35",
X"07D0",
X"0000",
X"F830",
X"F254",
X"F060",
X"F254",
X"F7B3",
X"FE89",
X"04E2",
X"08CA",
X"09C4",
X"07D0",
X"03E8",
X"FF83",
X"FC18",
X"FA24",
X"F9A7",
X"FAA1",
X"FC18",
X"FD8F",
X"FF06",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"007D",
X"0271",
X"055F",
X"0947",
X"0BB8",
X"0C35",
X"08CA",
X"01F4",
X"FA24",
X"F3CB",
X"F0DD",
X"F254",
X"F6B9",
X"FD8F",
X"03E8",
X"084D",
X"0947",
X"07D0",
X"0465",
X"0000",
X"FC18",
X"FA24",
X"F92A",
X"FA24",
X"FB9B",
X"FD8F",
X"FF83",
X"007D",
X"0177",
X"0177",
X"00FA",
X"007D",
X"007D",
X"01F4",
X"0465",
X"07D0",
X"0A41",
X"0ABE",
X"07D0",
X"0271",
X"FC18",
X"F63C",
X"F2D1",
X"F34E",
X"F736",
X"FC95",
X"02EE",
X"06D6",
X"084D",
X"0753",
X"03E8",
X"0000",
X"FC95",
X"FA24",
X"F92A",
X"FA24",
X"FB9B",
X"FD8F",
X"FF83",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0177",
X"03E8",
X"06D6",
X"09C4",
X"0A41",
X"084D",
X"036B",
X"FD8F",
X"F7B3",
X"F448",
X"F3CB",
X"F6B9",
X"FC18",
X"0177",
X"05DC",
X"0753",
X"06D6",
X"0465",
X"007D",
X"FD12",
X"FAA1",
X"F9A7",
X"FA24",
X"FB9B",
X"FD8F",
X"FF06",
X"007D",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"0177",
X"03E8",
X"0659",
X"08CA",
X"09C4",
X"07D0",
X"036B",
X"FE0C",
X"F8AD",
X"F542",
X"F448",
X"F63C",
X"FB1E",
X"007D",
X"04E2",
X"0753",
X"06D6",
X"0465",
X"00FA",
X"FD8F",
X"FB1E",
X"FA24",
X"FAA1",
X"FB9B",
X"FD8F",
X"FF83",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0177",
X"03E8",
X"06D6",
X"0947",
X"0947",
X"0753",
X"02EE",
X"FD8F",
X"F8AD",
X"F542",
X"F448",
X"F6B9",
X"FB1E",
X"007D",
X"04E2",
X"06D6",
X"06D6",
X"0465",
X"007D",
X"FD12",
X"FAA1",
X"F9A7",
X"FAA1",
X"FC18",
X"FE0C",
X"0000",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"007D",
X"01F4",
X"03E8",
X"06D6",
X"08CA",
X"0947",
X"06D6",
X"01F4",
X"FC95",
X"F830",
X"F542",
X"F542",
X"F7B3",
X"FC18",
X"0177",
X"055F",
X"06D6",
X"0659",
X"03E8",
X"007D",
X"FC95",
X"FAA1",
X"F9A7",
X"FAA1",
X"FC95",
X"FE0C",
X"0000",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"0177",
X"0271",
X"0465",
X"06D6",
X"084D",
X"07D0",
X"04E2",
X"007D",
X"FB9B",
X"F7B3",
X"F5BF",
X"F63C",
X"F92A",
X"FD8F",
X"01F4",
X"055F",
X"06D6",
X"05DC",
X"036B",
X"0000",
X"FC95",
X"FAA1",
X"FA24",
X"FAA1",
X"FC18",
X"FE0C",
X"FF83",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"01F4",
X"036B",
X"055F",
X"06D6",
X"07D0",
X"06D6",
X"036B",
X"FE89",
X"F9A7",
X"F6B9",
X"F5BF",
X"F736",
X"FAA1",
X"FF06",
X"036B",
X"05DC",
X"0659",
X"055F",
X"02EE",
X"FF83",
X"FC95",
X"FAA1",
X"FAA1",
X"FB1E",
X"FC95",
X"FE89",
X"0000",
X"00FA",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"02EE",
X"03E8",
X"055F",
X"0659",
X"0659",
X"0465",
X"00FA",
X"FC95",
X"F8AD",
X"F6B9",
X"F736",
X"F92A",
X"FC95",
X"00FA",
X"0465",
X"05DC",
X"0659",
X"0465",
X"01F4",
X"FE89",
X"FC18",
X"FAA1",
X"FAA1",
X"FB9B",
X"FD12",
X"FE89",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"03E8",
X"04E2",
X"05DC",
X"0659",
X"055F",
X"0271",
X"FE0C",
X"FA24",
X"F736",
X"F6B9",
X"F830",
X"FB1E",
X"FF06",
X"02EE",
X"05DC",
X"0659",
X"05DC",
X"03E8",
X"00FA",
X"FE0C",
X"FC18",
X"FB1E",
X"FAA1",
X"FB9B",
X"FD12",
X"FE89",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"0465",
X"04E2",
X"05DC",
X"05DC",
X"04E2",
X"01F4",
X"FE89",
X"FAA1",
X"F7B3",
X"F6B9",
X"F7B3",
X"FAA1",
X"FE0C",
X"01F4",
X"04E2",
X"0659",
X"0659",
X"04E2",
X"0271",
X"FF83",
X"FD12",
X"FB9B",
X"FB1E",
X"FB1E",
X"FC18",
X"FD12",
X"FE89",
X"0000",
X"0177",
X"02EE",
X"03E8",
X"04E2",
X"0659",
X"06D6",
X"06D6",
X"04E2",
X"01F4",
X"FD8F",
X"F92A",
X"F6B9",
X"F63C",
X"F7B3",
X"FAA1",
X"FE89",
X"01F4",
X"04E2",
X"0659",
X"0659",
X"055F",
X"036B",
X"00FA",
X"FE89",
X"FC95",
X"FB9B",
X"FB1E",
X"FB1E",
X"FC18",
X"FD8F",
X"FF83",
X"00FA",
X"02EE",
X"0465",
X"0659",
X"0753",
X"07D0",
X"06D6",
X"0465",
X"007D",
X"FC18",
X"F830",
X"F5BF",
X"F5BF",
X"F7B3",
X"FB1E",
X"FF06",
X"02EE",
X"055F",
X"06D6",
X"06D6",
X"05DC",
X"036B",
X"00FA",
X"FF06",
X"FD12",
X"FB9B",
X"FB1E",
X"FB1E",
X"FC18",
X"FD8F",
X"FF06",
X"007D",
X"0271",
X"0465",
X"0659",
X"07D0",
X"084D",
X"0753",
X"03E8",
X"FF83",
X"FAA1",
X"F736",
X"F542",
X"F5BF",
X"F830",
X"FB9B",
X"FF83",
X"0271",
X"04E2",
X"06D6",
X"06D6",
X"05DC",
X"03E8",
X"0177",
X"FF83",
X"FE0C",
X"FC95",
X"FB9B",
X"FB1E",
X"FB9B",
X"FC95",
X"FE0C",
X"0000",
X"01F4",
X"03E8",
X"05DC",
X"07D0",
X"08CA",
X"07D0",
X"04E2",
X"007D",
X"FB1E",
X"F736",
X"F542",
X"F5BF",
X"F7B3",
X"FAA1",
X"FE89",
X"01F4",
X"04E2",
X"0659",
X"0659",
X"05DC",
X"03E8",
X"01F4",
X"0000",
X"FE89",
X"FD12",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FD8F",
X"FE89",
X"007D",
X"02EE",
X"055F",
X"07D0",
X"0947",
X"08CA",
X"0659",
X"01F4",
X"FC18",
X"F7B3",
X"F4C5",
X"F4C5",
X"F63C",
X"F9A7",
X"FD8F",
X"00FA",
X"0465",
X"0659",
X"06D6",
X"05DC",
X"0465",
X"02EE",
X"00FA",
X"FF83",
X"FE0C",
X"FC95",
X"FC18",
X"FB9B",
X"FC18",
X"FD12",
X"FE89",
X"007D",
X"0271",
X"04E2",
X"06D6",
X"08CA",
X"08CA",
X"0753",
X"036B",
X"FE0C",
X"F92A",
X"F5BF",
X"F4C5",
X"F542",
X"F830",
X"FB9B",
X"0000",
X"036B",
X"05DC",
X"06D6",
X"0659",
X"04E2",
X"036B",
X"0177",
X"0000",
X"FE89",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FD12",
X"FE0C",
X"FF83",
X"00FA",
X"03E8",
X"0659",
X"08CA",
X"09C4",
X"08CA",
X"055F",
X"FF83",
X"F9A7",
X"F542",
X"F34E",
X"F448",
X"F6B9",
X"FAA1",
X"FF83",
X"036B",
X"05DC",
X"06D6",
X"0659",
X"055F",
X"036B",
X"01F4",
X"0000",
X"FF06",
X"FE0C",
X"FD12",
X"FC95",
X"FC18",
X"FC95",
X"FD8F",
X"FF06",
X"00FA",
X"036B",
X"0659",
X"08CA",
X"09C4",
X"08CA",
X"055F",
X"FF83",
X"F9A7",
X"F5BF",
X"F3CB",
X"F448",
X"F6B9",
X"FAA1",
X"FF06",
X"02EE",
X"055F",
X"0659",
X"0659",
X"04E2",
X"036B",
X"01F4",
X"007D",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE89",
X"007D",
X"02EE",
X"055F",
X"07D0",
X"0947",
X"08CA",
X"055F",
X"007D",
X"FAA1",
X"F63C",
X"F448",
X"F448",
X"F63C",
X"FA24",
X"FE89",
X"0271",
X"04E2",
X"0659",
X"05DC",
X"04E2",
X"036B",
X"01F4",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FE0C",
X"0000",
X"01F4",
X"0465",
X"06D6",
X"08CA",
X"0947",
X"0753",
X"02EE",
X"FD8F",
X"F830",
X"F542",
X"F448",
X"F542",
X"F830",
X"FC95",
X"00FA",
X"0465",
X"0659",
X"0659",
X"055F",
X"036B",
X"01F4",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FD8F",
X"FE89",
X"007D",
X"036B",
X"05DC",
X"07D0",
X"0947",
X"08CA",
X"05DC",
X"00FA",
X"FB9B",
X"F736",
X"F4C5",
X"F4C5",
X"F6B9",
X"FA24",
X"FE0C",
X"01F4",
X"04E2",
X"05DC",
X"055F",
X"0465",
X"0271",
X"00FA",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FF06",
X"00FA",
X"036B",
X"05DC",
X"084D",
X"0947",
X"084D",
X"0465",
X"FF06",
X"FA24",
X"F6B9",
X"F542",
X"F5BF",
X"F830",
X"FB9B",
X"0000",
X"036B",
X"055F",
X"05DC",
X"04E2",
X"036B",
X"0177",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE89",
X"0000",
X"01F4",
X"04E2",
X"0753",
X"08CA",
X"08CA",
X"0659",
X"01F4",
X"FC95",
X"F830",
X"F5BF",
X"F4C5",
X"F6B9",
X"FA24",
X"FE0C",
X"01F4",
X"04E2",
X"05DC",
X"055F",
X"03E8",
X"01F4",
X"007D",
X"FF06",
X"FE89",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF83",
X"0177",
X"03E8",
X"0659",
X"084D",
X"08CA",
X"06D6",
X"036B",
X"FE89",
X"F9A7",
X"F63C",
X"F542",
X"F63C",
X"F8AD",
X"FC95",
X"007D",
X"036B",
X"055F",
X"05DC",
X"0465",
X"02EE",
X"00FA",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE89",
X"0000",
X"0271",
X"04E2",
X"06D6",
X"084D",
X"07D0",
X"055F",
X"0177",
X"FD12",
X"F92A",
X"F6B9",
X"F63C",
X"F7B3",
X"FAA1",
X"FE0C",
X"0177",
X"03E8",
X"055F",
X"04E2",
X"036B",
X"01F4",
X"007D",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF83",
X"00FA",
X"0271",
X"04E2",
X"06D6",
X"07D0",
X"0753",
X"04E2",
X"0177",
X"FD8F",
X"F9A7",
X"F736",
X"F63C",
X"F7B3",
X"FAA1",
X"FE0C",
X"0177",
X"03E8",
X"055F",
X"04E2",
X"036B",
X"0177",
X"FF83",
X"FE0C",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"007D",
X"0271",
X"04E2",
X"06D6",
X"07D0",
X"0753",
X"055F",
X"01F4",
X"FD8F",
X"F9A7",
X"F6B9",
X"F63C",
X"F7B3",
X"FAA1",
X"FE89",
X"01F4",
X"0465",
X"055F",
X"04E2",
X"02EE",
X"00FA",
X"FF06",
X"FE0C",
X"FD8F",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"0000",
X"0271",
X"04E2",
X"0753",
X"084D",
X"084D",
X"05DC",
X"01F4",
X"FD8F",
X"F8AD",
X"F5BF",
X"F542",
X"F736",
X"FB1E",
X"FF83",
X"02EE",
X"055F",
X"05DC",
X"04E2",
X"02EE",
X"007D",
X"FF06",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FF06",
X"007D",
X"02EE",
X"055F",
X"07D0",
X"08CA",
X"07D0",
X"055F",
X"00FA",
X"FC18",
X"F7B3",
X"F542",
X"F542",
X"F7B3",
X"FB9B",
X"0000",
X"036B",
X"055F",
X"055F",
X"0465",
X"0271",
X"007D",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FF83",
X"00FA",
X"036B",
X"05DC",
X"07D0",
X"08CA",
X"07D0",
X"0465",
X"FF83",
X"FAA1",
X"F6B9",
X"F542",
X"F5BF",
X"F830",
X"FC18",
X"0000",
X"036B",
X"055F",
X"05DC",
X"04E2",
X"02EE",
X"0177",
X"0000",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FE0C",
X"FE89",
X"0000",
X"0271",
X"04E2",
X"06D6",
X"084D",
X"084D",
X"06D6",
X"036B",
X"FE89",
X"FA24",
X"F6B9",
X"F542",
X"F63C",
X"F8AD",
X"FC95",
X"007D",
X"03E8",
X"055F",
X"055F",
X"0465",
X"0271",
X"007D",
X"FF06",
X"FE0C",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"007D",
X"01F4",
X"0465",
X"0659",
X"07D0",
X"084D",
X"0659",
X"0271",
X"FE0C",
X"FA24",
X"F736",
X"F5BF",
X"F6B9",
X"F92A",
X"FD12",
X"007D",
X"036B",
X"055F",
X"055F",
X"03E8",
X"01F4",
X"0000",
X"FF06",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"0000",
X"0271",
X"04E2",
X"0753",
X"08CA",
X"08CA",
X"06D6",
X"036B",
X"FE89",
X"FA24",
X"F6B9",
X"F542",
X"F63C",
X"F92A",
X"FD12",
X"00FA",
X"0465",
X"05DC",
X"055F",
X"03E8",
X"01F4",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE89",
X"0000",
X"01F4",
X"04E2",
X"06D6",
X"084D",
X"084D",
X"06D6",
X"036B",
X"FE89",
X"F9A7",
X"F63C",
X"F4C5",
X"F63C",
X"F9A7",
X"FD8F",
X"0177",
X"0465",
X"05DC",
X"055F",
X"03E8",
X"01F4",
X"0000",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FF06",
X"00FA",
X"02EE",
X"05DC",
X"07D0",
X"08CA",
X"084D",
X"05DC",
X"01F4",
X"FD12",
X"F8AD",
X"F542",
X"F4C5",
X"F6B9",
X"FA24",
X"FE89",
X"0271",
X"055F",
X"05DC",
X"055F",
X"03E8",
X"01F4",
X"0000",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FF06",
X"00FA",
X"036B",
X"05DC",
X"07D0",
X"0947",
X"08CA",
X"05DC",
X"00FA",
X"FB9B",
X"F6B9",
X"F4C5",
X"F4C5",
X"F736",
X"FB1E",
X"FF83",
X"036B",
X"05DC",
X"0659",
X"055F",
X"036B",
X"0177",
X"FF83",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"0000",
X"0177",
X"03E8",
X"0659",
X"07D0",
X"08CA",
X"07D0",
X"04E2",
X"007D",
X"FB1E",
X"F736",
X"F542",
X"F542",
X"F7B3",
X"FB9B",
X"0000",
X"036B",
X"05DC",
X"0659",
X"05DC",
X"03E8",
X"0177",
X"FF83",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"0000",
X"01F4",
X"0465",
X"0659",
X"084D",
X"08CA",
X"07D0",
X"0465",
X"0000",
X"FB1E",
X"F736",
X"F5BF",
X"F63C",
X"F8AD",
X"FC95",
X"007D",
X"036B",
X"05DC",
X"05DC",
X"04E2",
X"02EE",
X"00FA",
X"FF06",
X"FE0C",
X"FD8F",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FF06",
X"007D",
X"01F4",
X"0465",
X"0659",
X"07D0",
X"08CA",
X"0753",
X"03E8",
X"FF06",
X"F9A7",
X"F6B9",
X"F5BF",
X"F6B9",
X"F9A7",
X"FD12",
X"0177",
X"0465",
X"0659",
X"0659",
X"04E2",
X"02EE",
X"007D",
X"FF06",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE0C",
X"FF06",
X"FF83",
X"00FA",
X"0271",
X"0465",
X"0659",
X"0753",
X"0753",
X"0659",
X"02EE",
X"FE89",
X"FA24",
X"F736",
X"F6B9",
X"F7B3",
X"FA24",
X"FD8F",
X"00FA",
X"03E8",
X"055F",
X"055F",
X"03E8",
X"01F4",
X"0000",
X"FE0C",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"0271",
X"03E8",
X"05DC",
X"06D6",
X"0753",
X"0659",
X"02EE",
X"FE89",
X"FA24",
X"F6B9",
X"F5BF",
X"F736",
X"FA24",
X"FE0C",
X"01F4",
X"04E2",
X"0659",
X"05DC",
X"0465",
X"01F4",
X"0000",
X"FE0C",
X"FD12",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"0271",
X"036B",
X"04E2",
X"05DC",
X"05DC",
X"04E2",
X"01F4",
X"FE89",
X"FB1E",
X"F8AD",
X"F7B3",
X"F8AD",
X"FB1E",
X"FE89",
X"0177",
X"0465",
X"055F",
X"055F",
X"03E8",
X"01F4",
X"FF83",
X"FE0C",
X"FD12",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"02EE",
X"0465",
X"055F",
X"055F",
X"0465",
X"0271",
X"FF83",
X"FC95",
X"FA24",
X"F8AD",
X"F9A7",
X"FB9B",
X"FE89",
X"0177",
X"036B",
X"04E2",
X"0465",
X"036B",
X"0177",
X"FF83",
X"FE0C",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"02EE",
X"03E8",
X"04E2",
X"04E2",
X"03E8",
X"0177",
X"FE89",
X"FC18",
X"FA24",
X"F9A7",
X"FA24",
X"FC95",
X"FF83",
X"01F4",
X"03E8",
X"04E2",
X"0465",
X"02EE",
X"00FA",
X"FF06",
X"FD8F",
X"FC95",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"036B",
X"0271",
X"007D",
X"FE89",
X"FC95",
X"FB1E",
X"FAA1",
X"FB9B",
X"FD8F",
X"0000",
X"01F4",
X"036B",
X"03E8",
X"036B",
X"01F4",
X"007D",
X"FF06",
X"FD8F",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"036B",
X"02EE",
X"0177",
X"FF83",
X"FD12",
X"FB9B",
X"FB1E",
X"FB1E",
X"FC95",
X"FE89",
X"00FA",
X"02EE",
X"0465",
X"0465",
X"036B",
X"01F4",
X"0000",
X"FE89",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"00FA",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"00FA",
X"FF83",
X"FE0C",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FE0C",
X"0000",
X"01F4",
X"036B",
X"03E8",
X"03E8",
X"02EE",
X"0177",
X"FF83",
X"FE0C",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE89",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"0177",
X"007D",
X"FF06",
X"FD8F",
X"FC95",
X"FC18",
X"FC95",
X"FD8F",
X"FF06",
X"00FA",
X"0271",
X"036B",
X"03E8",
X"036B",
X"01F4",
X"007D",
X"FF06",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"007D",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0271",
X"01F4",
X"00FA",
X"FF83",
X"FE0C",
X"FD12",
X"FC18",
X"FC18",
X"FD12",
X"FE89",
X"007D",
X"01F4",
X"036B",
X"03E8",
X"036B",
X"0271",
X"00FA",
X"FF83",
X"FE0C",
X"FD12",
X"FD12",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"0177",
X"007D",
X"FF06",
X"FD8F",
X"FC18",
X"FB9B",
X"FC18",
X"FD8F",
X"FF06",
X"00FA",
X"02EE",
X"03E8",
X"03E8",
X"02EE",
X"01F4",
X"0000",
X"FE89",
X"FD8F",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"00FA",
X"FF83",
X"FE0C",
X"FD12",
X"FC18",
X"FC18",
X"FC95",
X"FE0C",
X"0000",
X"01F4",
X"036B",
X"03E8",
X"03E8",
X"02EE",
X"0177",
X"FF83",
X"FE0C",
X"FD12",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"007D",
X"FF06",
X"FE0C",
X"FD12",
X"FC95",
X"FC95",
X"FD8F",
X"FF06",
X"007D",
X"0271",
X"036B",
X"036B",
X"036B",
X"0271",
X"00FA",
X"FF83",
X"FE0C",
X"FD12",
X"FD12",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FD8F",
X"FF06",
X"007D",
X"01F4",
X"02EE",
X"036B",
X"036B",
X"0271",
X"0177",
X"0000",
X"FE89",
X"FD8F",
X"FD12",
X"FD12",
X"FD8F",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"01F4",
X"0271",
X"01F4",
X"01F4",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"0177",
X"0271",
X"02EE",
X"036B",
X"02EE",
X"01F4",
X"007D",
X"FF83",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FE0C",
X"FF06",
X"007D",
X"0177",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FD8F",
X"FE0C",
X"FF83",
X"007D",
X"0177",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE0C",
X"FD8F",
X"FD12",
X"FD8F",
X"FE89",
X"0000",
X"00FA",
X"01F4",
X"0271",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83"


 );

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
--      if (ENA='1') then
		Q_tmp <= sin_table(conv_integer(ADDR));
--      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end arch;