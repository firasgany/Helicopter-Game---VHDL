library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;
-- Alex Grinshpun July 24 2017 
-- Dudy Nov 13 2017


entity cieling_draw is
port 	(
		
	   CLK      : in std_logic;
		RESETn	: in std_logic;
		oCoord_X : in integer;
		oCoord_Y : in integer;
		drawing_request : out std_logic ;
		mVGA_RGB	: out std_logic_vector(7 downto 0) --	,//	VGA composite RGB
	);
end cieling_draw;

architecture behav of cieling_draw is 

-- Constants for frame drawing
--constant	x_frame	: integer :=	639;
--constant	y_frame	: integer :=	479;
----constant	int_frame	: integer :=	10;

signal mVGA_R	: std_logic_vector(2 downto 0); --	,	 			//	VGA Red[2:0]
signal mVGA_G	: std_logic_vector(2 downto 0); --	,	 			//	VGA Green[2:0]
signal mVGA_B	: std_logic_vector(1 downto 0); --	,  			//	VGA Blue[1:0]


	
begin
mVGA_RGB <=  mVGA_R & mVGA_G &  mVGA_B ;

process (RESETn, CLK, oCoord_X,oCoord_Y)

type RAM_ARRAY is array (0 to 15981) of integer range 0 to 100;
constant height_value : RAM_ARRAY := (

46,46,44,43,42,43,44,46,46,46,46,46,46,46,46,46,46,46,46,46,46,46,44,43,42,42,42,42,42,42,42,42,42,42,42,42,42,42,42,42,42,42,42,42,42,42,42,42,42,42,42,43,44,47,48,51,52,54,54,54,54,54,54,54,54,54,54,54,55,56,58,58,58,58,56,56,56,58,58,58,56,55,52,51,50,50,50,50,50,50,50,50,50,48,47,46,46,46,46,46,44,43,42,42,42,42,42,42,42,42,42,42,40,39,39,40,42,43,44,44,42,40,39,39,38,38,38,38,38,38,38,38,38,36,35,34,34,34,34,34,34,32,31,30,30,30,28,27,27,28,28,27,26,26,27,28,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,31,32,34,32,31,31,32,34,34,34,34,32,31,31,32,34,34,34,34,34,35,35,34,32,32,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,32,31,30,30,28,28,28,30,30,30,30,30,28,28,28,31,32,34,34,32,31,30,28,28,27,27,24,23,22,23,24,24,23,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,23,23,23,22,22,22,23,24,26,26,26,26,26,27,28,30,30,30,30,30,31,32,34,32,31,30,30,30,28,27,26,26,26,24,23,22,22,22,22,22,22,22,23,24,26,26,24,22,20,20,23,24,26,26,26,26,26,26,26,24,22,19,18,18,18,18,19,20,23,24,26,26,26,26,26,26,26,26,26,26,26,24,23,22,20,19,18,18,18,18,18,18,18,16,16,16,18,18,18,18,18,18,18,16,15,14,12,11,10,10,10,10,10,10,10,10,10,10,10,10,8,7,6,7,8,8,7,6,4,3,2,3,4,6,6,6,4,3,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,4,4,5,6,8,9,10,12,12,12,12,12,12,12,12,12,12,12,12,10,9,6,5,4,4,5,6,8,8,8,8,8,8,8,8,8,8,8,8,6,5,4,4,4,4,5,6,8,8,8,8,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,6,8,8,6,5,4,4,4,3,3,3,5,6,8,8,8,8,8,8,8,8,8,8,8,9,12,14,16,16,16,16,16,16,16,16,16,16,16,17,18,20,21,24,28,30,32,32,32,30,28,25,24,24,24,24,25,26,26,25,22,21,20,20,18,18,20,22,24,24,24,24,24,24,24,24,24,22,22,22,24,24,24,25,26,28,26,25,24,24,24,24,22,21,20,20,20,20,18,17,16,16,16,16,16,16,16,16,16,16,16,16,17,18,20,20,20,20,20,20,20,20,18,17,16,16,16,16,16,16,16,16,16,16,16,16,14,13,12,12,12,10,9,9,12,14,17,18,20,18,17,16,16,16,16,16,14,13,10,8,5,4,4,3,3,3,4,4,4,5,6,8,8,8,8,8,8,8,8,8,8,8,9,10,12,12,12,12,12,12,12,12,10,9,9,10,12,12,13,14,16,16,14,13,13,14,16,16,16,16,16,17,20,22,24,24,24,24,24,24,24,24,25,26,28,28,28,28,28,29,30,32,30,29,28,28,29,29,29,28,29,30,32,32,33,34,36,36,36,36,37,38,40,40,40,41,42,44,44,45,46,48,48,48,48,48,46,45,44,44,44,44,44,45,46,48,48,48,48,48,46,45,45,45,45,44,44,44,44,44,44,44,44,45,46,48,48,48,48,48,46,46,46,48,48,49,50,52,52,52,52,52,52,52,52,52,52,52,52,52,52,52,53,54,56,56,56,56,56,56,56,57,57,57,57,58,60,60,60,60,60,60,60,61,62,64,64,64,64,64,64,64,64,64,64,65,66,68,68,68,68,66,65,65,66,68,68,66,65,64,64,64,64,64,64,64,64,62,61,58,57,56,56,56,56,56,54,53,52,50,49,48,48,48,48,48,48,48,49,50,53,54,56,56,56,56,54,52,49,48,48,48,49,50,52,50,50,50,53,56,58,60,60,60,60,60,58,57,56,56,56,56,56,56,56,57,58,60,60,60,60,60,60,60,60,60,60,60,60,61,62,64,64,64,64,65,66,68,68,68,66,65,64,64,64,64,65,66,66,65,64,64,64,64,64,64,64,64,64,65,66,68,68,68,69,70,72,72,72,72,73,74,76,77,80,82,84,84,84,84,85,86,88,88,88,86,85,82,81,80,80,80,80,80,80,80,80,80,80,80,80,80,80,78,77,76,76,76,76,76,76,76,76,76,74,73,70,69,68,68,66,66,66,68,68,68,68,68,68,68,68,68,68,68,68,68,68,66,65,64,64,64,64,64,64,64,64,65,66,68,68,68,68,68,68,68,68,68,68,68,68,68,66,65,64,64,62,61,60,60,60,60,60,60,58,57,56,56,56,56,56,56,56,56,57,58,60,61,62,62,61,60,61,62,64,65,66,68,68,68,68,66,65,64,64,65,66,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,66,66,66,68,68,68,68,68,69,70,72,72,72,72,72,72,72,72,72,73,74,76,76,74,72,68,65,64,64,64,64,64,64,62,60,57,56,57,58,60,61,62,64,64,64,64,64,64,64,62,62,62,65,65,65,64,64,64,62,61,60,61,64,66,68,66,65,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,65,66,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,66,65,64,62,61,60,60,60,60,60,60,60,60,60,61,62,64,64,64,62,61,60,60,60,60,60,60,58,57,56,56,56,56,56,56,56,54,53,52,52,52,52,52,52,53,54,56,56,57,58,60,58,57,56,56,56,56,56,56,56,56,56,56,56,56,56,56,57,58,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,58,57,56,57,57,56,53,52,52,52,52,53,54,56,56,56,54,53,52,52,50,49,48,48,48,49,52,56,60,62,64,64,64,65,66,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,66,64,61,60,60,58,58,58,58,57,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,57,57,57,57,58,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,58,57,56,56,56,54,53,52,52,52,53,54,56,56,56,56,56,56,56,56,56,56,56,54,53,52,50,49,46,45,44,44,44,44,44,42,41,40,40,40,40,40,40,40,40,40,40,40,40,40,40,41,44,46,48,49,50,52,50,49,49,50,52,52,52,52,52,52,50,49,48,48,48,48,48,49,50,52,52,52,52,50,50,49,49,46,45,44,44,44,45,46,48,48,48,48,48,48,48,48,48,48,49,50,52,52,52,52,52,52,52,52,53,54,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,57,58,60,60,60,61,62,64,65,66,68,68,68,68,68,66,65,65,66,68,68,68,68,68,68,68,68,66,65,64,64,64,64,62,61,60,60,60,60,60,60,61,62,64,64,64,64,64,64,62,61,60,61,61,61,61,61,61,60,60,60,60,60,60,60,58,57,56,54,53,52,52,52,52,52,52,52,53,54,56,56,56,56,56,56,56,56,54,53,53,54,54,54,54,56,56,56,56,56,56,56,54,53,50,50,50,52,52,52,52,52,50,49,48,48,48,48,48,48,48,46,45,44,44,44,44,42,41,40,40,40,40,40,40,40,38,36,33,32,32,32,32,32,30,29,28,28,28,26,25,24,24,24,24,22,21,20,20,20,20,20,20,20,18,17,16,16,16,17,18,21,22,24,24,24,24,25,26,28,28,28,28,26,24,21,20,20,20,20,20,20,20,20,20,20,20,20,21,22,24,24,24,24,24,24,24,24,24,24,24,24,22,22,22,24,24,24,24,24,25,26,28,28,28,28,28,28,28,28,28,28,29,30,32,32,33,34,36,36,36,36,37,38,40,40,38,37,36,36,36,36,36,36,36,37,38,40,38,37,37,38,40,40,40,40,40,40,40,40,40,40,41,42,44,45,46,49,50,52,53,54,56,56,57,58,61,62,62,61,60,60,60,60,60,58,57,56,57,58,60,60,60,60,60,60,60,60,60,60,60,60,60,58,57,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,57,60,62,64,64,64,64,64,62,61,60,60,60,60,60,58,58,58,60,60,60,60,58,57,56,56,56,56,56,56,54,53,52,52,52,52,52,53,54,56,56,54,53,52,52,52,52,52,52,52,53,54,56,56,56,56,56,56,56,56,56,56,56,56,56,57,60,62,64,64,64,64,64,64,64,64,64,64,62,61,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,61,62,64,64,62,61,60,60,60,60,60,60,60,60,60,60,60,60,60,61,62,65,66,68,68,68,68,68,68,68,69,69,70,70,72,72,72,72,72,72,72,72,72,72,72,72,72,72,72,72,72,72,70,69,68,68,68,68,68,68,68,68,68,68,69,70,72,72,70,68,65,64,62,62,62,62,61,61,62,62,61,60,60,60,60,60,60,60,60,61,62,64,64,64,64,64,64,64,64,64,64,64,64,62,61,60,60,60,58,57,56,56,54,53,52,52,52,52,52,52,52,52,52,52,53,54,56,56,56,56,56,56,56,57,58,60,60,58,56,53,52,52,52,52,52,52,52,52,52,52,52,52,52,52,53,54,56,57,57,57,56,56,56,56,56,57,58,61,64,66,68,68,66,65,64,64,64,65,66,68,68,68,68,68,68,68,68,68,69,70,73,73,74,74,76,76,76,76,76,76,76,76,76,76,74,73,72,72,70,69,68,68,69,70,73,74,76,76,76,76,76,76,76,76,76,74,73,72,72,72,70,69,68,68,68,68,68,68,68,69,70,70,69,68,69,70,70,69,68,68,68,69,70,72,72,72,73,74,76,76,76,74,73,72,72,72,72,72,72,70,69,68,68,68,69,70,72,72,72,72,72,70,69,66,65,64,64,64,64,65,68,70,72,72,72,72,72,72,72,72,73,74,76,76,76,76,77,78,80,80,80,80,80,80,80,80,80,80,80,80,80,80,80,80,80,80,80,80,78,77,76,76,76,76,76,76,76,76,76,76,76,77,78,80,78,77,76,76,77,78,80,80,80,80,78,77,74,73,73,76,78,80,80,80,81,82,84,84,85,86,88,88,88,88,89,90,92,92,93,96,98,100,100,98,97,96,96,96,96,96,96,96,96,97,98,100,98,97,96,96,97,98,100,100,100,100,100,100,100,100,98,97,96,94,94,94,96,96,96,96,96,96,96,96,96,96,96,96,96,96,94,93,90,89,86,85,84,84,84,84,84,84,84,84,84,84,84,84,82,82,82,84,84,84,84,84,84,84,84,84,84,84,84,84,84,85,86,88,86,85,84,84,84,84,84,85,86,88,88,88,88,89,90,92,93,94,96,96,94,93,92,92,92,92,92,92,92,92,92,92,90,89,88,88,88,89,90,92,93,94,94,92,90,89,88,85,84,82,81,80,80,80,80,80,78,76,73,72,72,72,72,72,70,69,68,68,68,68,69,72,73,72,69,68,66,65,64,64,64,64,64,62,61,58,57,56,56,56,56,56,56,56,56,56,54,54,54,56,56,56,56,56,57,58,60,58,57,56,56,56,56,56,54,53,52,53,54,56,56,56,56,56,54,52,49,48,48,48,48,48,46,44,41,40,38,37,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,37,38,40,40,40,40,40,40,40,40,40,40,40,40,40,40,38,37,36,36,34,34,34,36,34,33,30,28,26,26,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,26,25,24,25,26,28,26,25,24,22,21,20,20,20,20,21,22,24,24,24,24,24,24,24,24,24,22,21,20,20,20,20,20,20,21,22,24,24,24,24,24,24,24,24,24,22,21,20,20,20,20,20,21,22,24,24,24,22,21,20,21,22,25,26,28,28,26,25,24,24,24,24,24,24,24,24,24,24,24,24,24,25,26,28,28,26,25,24,24,24,22,21,20,20,20,20,20,20,20,20,20,20,21,21,21,20,20,20,20,20,20,18,16,13,10,9,8,8,8,9,10,10,9,8,8,9,10,10,9,6,5,3,3,3,5,5,5,4,4,4,4,4,4,4,4,4,4,5,6,9,10,12,12,12,12,12,10,9,8,8,8,8,8,8,8,8,8,8,8,6,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,6,8,8,8,8,6,7,5,5,4,4,4,4,3,3,3,4,4,4,4,4,4,4,5,5,5,4,4,4,4,4,4,4,4,5,6,8,8,8,8,8,8,8,8,8,8,9,10,12,10,9,8,8,6,5,4,4,5,5,5,4,4,4,4,4,5,6,8,8,8,6,5,4,4,5,8,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,5,4,4,4,4,4,4,4,4,4,4,5,5,6,5,5,4,5,6,6,5,5,6,8,8,8,8,8,8,8,9,10,12,13,14,16,16,17,18,20,20,20,20,20,20,20,20,21,22,24,24,24,24,24,24,24,22,20,17,16,16,17,18,20,20,20,20,20,20,20,20,20,20,18,17,16,16,16,16,16,16,16,16,16,16,16,16,17,18,18,16,13,12,12,12,12,12,12,12,12,12,10,9,8,8,8,8,8,8,9,10,13,14,14,13,12,12,10,9,8,8,6,5,5,6,8,8,8,8,8,8,8,9,10,10,9,6,5,5,6,8,8,8,8,6,5,5,6,9,10,12,12,12,12,12,12,12,12,12,10,9,8,9,10,12,12,12,13,16,18,20,20,20,20,20,21,22,24,25,26,26,26,26,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,26,25,24,24,25,26,29,30,32,32,32,32,33,34,36,36,36,37,38,40,40,40,40,38,38,40,41,41,40,40,40,40,38,37,37,38,40,40,40,40,40,38,37,36,36,36,36,36,36,36,36,36,36,36,36,36,37,40,42,44,44,44,44,44,44,44,44,44,44,44,45,46,48,48,49,52,54,56,56,57,58,60,60,60,60,60,60,60,60,60,60,60,60,61,61,61,60,60,60,60,60,60,60,58,57,56,56,56,56,56,56,56,56,56,57,58,60,61,61,61,60,60,60,60,60,60,61,62,64,64,64,64,64,64,64,64,64,64,64,64,62,60,56,52,49,46,44,41,38,37,36,36,36,34,33,32,30,29,28,26,25,24,24,24,24,22,21,18,17,16,16,17,18,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,18,17,17,18,20,20,20,20,20,20,20,21,22,24,24,22,21,20,18,17,16,14,13,12,12,12,12,12,12,12,13,14,16,16,16,16,16,16,16,16,16,17,18,20,20,20,18,17,17,18,20,20,20,18,17,16,17,18,20,20,20,20,20,20,20,20,20,20,18,17,16,16,16,16,14,13,12,12,12,12,13,13,13,12,12,12,12,12,13,14,16,16,16,16,16,16,16,16,17,18,20,20,20,20,21,22,24,24,24,22,21,20,20,20,20,20,18,17,16,17,17,17,16,14,13,12,10,9,9,9,9,8,9,10,10,9,8,8,8,8,8,8,9,10,12,12,12,12,12,12,10,9,8,8,8,8,6,5,4,4,4,4,4,4,4,5,4,4,3,4,4,4,4,4,5,6,8,8,8,8,6,5,4,4,4,5,6,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,10,12,10,9,8,8,8,8,8,6,6,5,5,4,4,4,4,4,4,4,4,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,3,3,4,5,5,4,4,4,4,4,3,3,3,4,4,4,4,4,4,5,6,8,8,8,6,5,4,4,4,4,4,4,4,4,3,3,3,5,6,8,8,8,8,6,5,4,4,4,4,4,4,5,8,12,14,17,18,18,17,16,16,16,16,16,16,16,16,16,16,16,14,13,12,10,9,8,6,5,5,6,6,5,4,5,6,8,8,8,8,8,8,8,8,8,8,8,8,6,5,4,4,5,6,8,8,6,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,6,8,8,8,8,8,8,8,9,10,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,14,16,14,13,12,12,12,12,12,12,10,9,8,8,8,8,8,8,8,8,8,8,8,8,6,5,4,4,4,5,6,8,8,8,6,5,4,4,4,4,4,4,4,4,4,4,4,4,5,6,9,10,12,12,12,12,10,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,10,12,13,14,16,17,18,21,22,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,25,26,28,28,28,28,29,30,32,32,32,32,32,32,32,32,32,32,32,32,33,34,36,34,33,32,32,33,34,36,36,36,36,37,38,41,42,44,44,44,44,44,44,44,44,45,48,50,52,52,52,52,52,52,53,54,56,57,58,60,60,58,57,56,57,58,60,60,60,60,60,60,61,62,64,65,66,69,70,73,73,73,72,73,74,76,76,76,76,76,76,76,76,74,73,72,72,72,70,69,68,68,69,70,72,72,73,74,76,76,74,73,72,72,72,72,72,73,73,73,73,74,74,74,74,76,76,76,74,73,72,72,72,72,72,73,76,78,80,80,80,80,80,80,80,80,78,77,76,76,76,76,76,76,76,76,76,77,78,80,78,77,76,76,76,76,76,76,77,78,80,80,80,80,80,80,80,80,80,80,80,80,80,80,80,80,80,80,80,80,80,78,77,76,76,77,78,80,80,80,81,82,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,82,81,80,80,80,81,82,84,84,84,84,85,86,88,88,88,88,88,88,88,88,86,84,81,80,78,77,76,76,76,77,78,80,78,77,76,76,76,77,80,82,85,86,86,85,84,84,84,85,88,90,92,92,92,90,89,88,88,88,88,88,86,85,84,84,84,84,84,84,84,84,84,85,86,88,88,88,88,88,88,88,88,88,88,88,88,86,85,84,84,84,85,86,86,84,81,78,77,77,78,78,77,76,76,76,76,76,76,76,76,76,76,76,76,76,76,76,77,78,81,82,84,82,81,80,80,80,80,80,80,81,82,84,84,82,81,80,81,82,84,84,82,81,80,80,80,80,80,80,80,78,77,76,76,77,78,80,80,80,80,80,80,80,80,80,80,81,82,85,86,88,88,88,88,88,88,88,88,89,90,92,92,92,92,90,89,89,90,93,94,97,98,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,98,97,96,96,96,96,96,96,94,93,92,92,93,94,96,96,94,93,92,92,92,92,92,92,92,93,93,93,92,92,93,94,96,94,93,93,94,96,96,96,96,96,96,96,96,97,98,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,98,97,96,96,96,97,98,100,100,100,100,100,100,100,100,100,100,100,98,97,96,96,96,96,96,97,98,100,100,100,100,100,98,96,92,89,89,90,92,92,92,92,92,92,92,92,92,92,93,94,96,96,96,96,96,94,93,92,93,94,94,93,93,94,96,96,96,96,94,93,92,92,92,92,92,92,93,94,96,96,97,97,96,93,90,89,88,88,88,88,89,90,90,89,88,86,85,84,84,84,84,84,84,84,85,85,85,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,85,86,88,88,86,85,84,84,84,84,84,84,82,81,80,80,80,81,84,86,88,88,88,88,88,88,88,86,85,82,82,81,81,80,80,80,80,80,81,82,84,84,84,84,84,84,84,84,84,84,84,84,84,82,82,82,85,86,88,88,88,88,88,88,88,88,88,88,89,90,92,92,92,92,92,93,94,96,96,97,98,100,100,100,100,100,100,100,98,97,97,98,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,98,97,96,96,96,96,96,96,96,96,96,96,97,98,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,98,97,94,93,92,92,92,92,92,92,92,92,93,94,96,94,93,92,92,92,92,93,96,98,100,100,100,100,100,100,100,100,100,100,100,100,100,98,96,93,90,89,88,89,90,92,92,92,92,92,92,92,90,89,88,88,88,88,88,89,90,92,92,92,92,90,90,90,92,92,90,89,88,88,86,84,81,80,80,80,80,80,81,82,85,86,88,88,88,88,88,88,86,84,81,80,80,80,80,80,80,81,82,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,85,86,88,88,88,88,86,85,84,84,84,85,86,88,88,88,88,88,88,88,88,88,88,88,88,88,88,88,88,88,88,88,86,85,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,82,80,77,76,76,76,76,76,76,77,78,80,78,76,73,70,69,69,72,76,78,80,78,77,76,76,76,76,76,76,76,74,73,70,69,68,68,68,68,68,68,68,68,68,68,68,68,66,65,64,64,65,66,69,70,70,69,68,66,65,64,64,64,64,64,64,62,61,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,58,57,56,56,56,54,54,56,58,60,60,60,60,60,58,57,56,56,56,56,56,57,58,60,61,62,64,64,62,61,60,60,60,60,60,60,60,60,60,60,60,58,57,56,56,57,58,60,60,58,57,56,57,58,61,62,64,64,64,64,62,61,58,57,56,56,56,54,53,52,52,52,52,52,52,52,53,54,56,56,56,56,56,56,56,56,54,53,52,52,50,50,50,52,53,54,56,56,56,56,56,56,56,56,56,57,58,60,58,57,56,56,56,56,56,56,56,56,56,56,56,56,56,54,53,52,52,53,53,53,52,52,50,49,48,48,48,48,46,45,44,44,44,44,44,44,44,44,42,41,40,40,40,38,37,36,36,34,33,32,32,32,33,34,34,32,29,28,28,28,28,29,30,30,29,28,28,28,28,28,28,28,28,28,28,29,29,29,28,28,28,28,28,28,28,28,28,26,25,24,24,24,24,24,24,24,25,26,28,28,28,28,28,28,28,28,28,28,28,28,26,25,24,24,24,24,24,24,24,24,22,21,20,18,16,13,12,12,12,10,9,8,8,8,8,9,12,14,16,16,16,17,18,20,20,21,22,24,24,24,24,25,25,26,28,30,33,34,36,37,38,38,37,36,36,36,36,36,36,36,36,36,37,38,40,38,37,36,36,36,36,36,36,37,38,40,41,42,44,44,44,44,44,44,44,44,44,44,42,41,40,41,41,41,40,41,41,41,40,40,40,38,38,40,42,44,44,44,44,44,44,44,42,40,37,36,36,36,34,33,32,33,34,36,34,33,32,32,33,34,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,37,38,40,40,40,40,40,40,40,40,40,40,40,41,42,42,41,40,40,40,40,40,40,40,41,42,44,44,44,44,45,46,48,49,50,52,52,52,52,52,52,52,53,56,60,62,64,65,66,68,68,68,68,68,68,68,68,68,68,68,69,70,72,72,72,73,74,76,76,76,74,73,72,70,69,68,68,69,70,72,72,70,69,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,69,70,72,72,72,72,72,72,70,69,68,68,68,68,68,69,69,69,68,68,68,68,68,68,69,70,72,70,69,68,68,68,68,68,68,68,68,68,68,68,66,65,64,64,64,64,64,64,64,64,64,65,66,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,66,65,64,64,64,64,64,62,61,60,60,60,60,60,58,57,56,56,56,56,56,56,57,60,62,64,64,64,64,64,64,64,64,64,64,64,64,64,62,61,61,62,64,64,64,64,64,64,64,65,66,68,68,68,68,66,65,64,64,62,61,60,61,62,62,61,60,60,60,60,61,62,64,64,64,64,64,64,65,66,68,66,66,66,68,66,65,64,62,61,60,60,58,57,56,56,56,56,56,54,54,54,54,53,52,52,52,52,50,48,45,42,40,37,34,33,32,32,32,32,32,32,32,33,34,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,37,38,40,38,37,36,36,37,40,42,44,42,41,41,42,44,42,41,40,40,41,42,44,44,44,44,42,41,40,38,37,36,36,34,33,32,30,29,29,30,32,32,32,32,32,32,32,32,33,34,36,36,36,36,36,36,36,36,36,36,36,36,37,38,40,38,37,34,33,33,34,36,37,38,40,40,40,40,40,40,40,40,40,40,40,40,41,42,44,44,42,41,40,40,41,42,44,44,44,44,44,44,44,44,44,44,44,44,44,44,42,41,40,40,38,38,38,40,40,38,38,38,40,40,40,40,40,40,38,37,36,36,36,36,36,36,34,33,32,32,32,30,29,28,28,28,28,28,28,26,26,26,28,28,28,26,25,24,24,24,24,22,21,20,18,16,13,13,14,16,16,14,13,12,12,12,12,13,14,17,18,18,17,17,18,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,21,22,22,21,20,20,20,20,20,20,20,20,21,22,22,21,20,20,20,20,21,22,25,25,25,22,22,22,25,25,25,24,22,20,17,17,18,20,18,17,16,16,14,13,12,13,14,16,16,16,16,16,16,16,16,16,14,13,12,12,12,12,10,9,8,8,6,5,4,4,3,3,3,4,4,4,4,4,4,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,5,6,8,9,10,12,12,12,12,12,12,12,12,12,12,13,14,16,16,16,17,20,22,24,24,25,26,28,28,28,28,28,28,28,28,28,28,28,28,28,26,25,24,24,24,24,24,24,24,24,24,24,24,24,25,26,29,30,32,32,32,32,32,30,29,28,28,28,28,28,28,28,28,28,28,28,29,30,32,32,32,32,30,29,29,30,33,34,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,34,33,32,32,32,32,30,30,30,32,32,32,32,32,32,32,32,32,32,33,34,36,36,36,36,36,36,36,36,36,37,38,40,40,40,40,40,40,40,40,40,40,38,37,36,34,33,32,32,32,32,33,34,37,38,40,40,40,38,38,38,40,40,40,40,41,42,44,44,42,41,40,40,40,38,38,37,37,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,37,38,40,40,40,40,40,41,41,41,40,40,40,40,40,40,40,40,40,40,40,40,40,40,38,37,37,38,41,42,44,44,45,46,48,48,48,49,50,52,52,52,52,52,52,50,49,48,48,48,48,48,49,50,52,52,52,52,53,54,56,56,57,58,60,58,58,58,60,60,60,61,61,61,60,61,62,64,64,64,65,65,65,64,64,64,62,60,57,56,56,56,56,56,56,56,56,56,56,56,54,53,52,52,52,52,52,52,50,49,48,49,50,52,52,52,52,52,53,53,53,52,52,53,54,56,56,56,56,56,56,56,56,56,56,56,56,57,58,60,58,57,57,60,61,61,60,60,60,60,60,60,60,60,60,60,60,60,60,61,62,64,64,64,64,64,62,61,60,60,60,60,60,58,57,56,56,56,56,56,56,56,56,56,54,53,52,52,52,52,52,53,54,56,56,54,53,52,52,50,49,49,52,54,56,56,56,54,53,52,52,52,50,50,49,50,50,52,52,53,54,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,54,53,52,52,52,53,53,53,52,50,49,48,48,48,49,52,54,57,58,60,60,60,60,60,58,57,56,54,53,52,50,49,48,48,48,48,48,49,50,52,52,52,52,53,54,56,56,56,54,53,52,50,49,48,49,50,52,52,52,52,52,52,52,52,52,52,52,53,54,54,53,52,53,54,56,57,58,60,60,60,60,60,60,61,62,62,61,60,61,61,61,60,60,60,60,60,60,60,60,60,60,60,60,60,60,61,62,64,64,64,64,64,64,64,64,64,64,64,62,60,56,53,52,52,52,52,52,52,52,52,52,52,52,52,53,54,56,56,54,53,52,52,52,52,50,49,48,48,48,49,50,52,53,54,56,56,56,56,57,58,60,61,62,64,64,64,64,64,65,66,68,68,69,69,69,68,68,68,68,68,68,68,68,69,72,74,76,76,76,76,76,76,76,76,76,76,76,76,76,76,77,77,78,78,80,80,80,80,81,82,84,84,84,82,80,77,76,76,76,74,73,72,72,70,69,68,68,68,66,65,64,64,64,64,64,64,64,64,64,64,64,64,64,65,66,68,68,68,68,68,66,64,61,60,60,58,57,54,53,52,52,53,54,56,56,56,56,57,58,61,64,66,68,68,68,69,70,73,74,76,76,76,76,76,77,78,81,84,86,88,86,85,84,84,84,84,84,84,85,86,88,88,88,86,86,86,88,88,89,90,92,92,90,89,89,90,92,92,92,92,93,94,94,93,92,92,92,92,92,92,92,92,92,90,89,89,90,92,90,89,88,88,88,88,88,88,88,88,88,88,86,85,84,84,85,86,88,88,88,88,88,88,88,88,88,89,89,89,88,88,89,90,92,92,92,92,92,92,92,92,92,92,92,92,92,93,94,96,96,96,96,96,96,96,96,96,96,97,98,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,98,97,96,96,96,96,96,96,96,94,93,90,89,88,89,90,92,93,94,96,96,96,96,96,96,96,96,96,96,96,96,96,97,98,100,100,100,100,100,100,100,100,100,100,100,100,100,98,97,96,94,92,89,86,85,82,81,80,80,81,82,84,82,81,80,80,80,80,80,80,80,80,78,77,76,76,76,77,78,81,82,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,85,86,88,89,90,93,94,96,96,94,93,92,92,92,90,89,86,85,84,84,84,84,84,84,82,81,80,80,80,80,80,80,80,81,84,85,85,84,84,84,84,84,84,84,84,84,84,84,85,86,88,88,88,88,88,88,88,88,88,86,86,86,88,86,85,84,84,84,82,81,80,80,80,81,82,84,84,85,86,88,88,88,86,85,84,84,84,82,81,78,77,76,74,73,72,72,72,72,72,72,72,72,72,72,70,69,68,68,68,68,69,70,72,72,73,74,76,76,77,78,80,80,80,80,80,80,80,80,80,80,80,80,78,77,76,76,76,76,76,76,76,74,73,72,72,72,73,74,76,76,76,76,76,76,76,76,76,77,78,80,80,80,80,80,80,80,80,80,81,82,84,85,86,88,89,90,92,92,92,92,92,93,94,96,96,96,96,97,98,100,100,98,97,96,96,94,93,92,92,92,92,92,90,90,89,89,86,84,81,81,82,84,85,86,88,88,88,86,85,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,82,81,80,80,78,78,78,80,81,82,84,84,84,84,84,84,84,82,81,78,77,76,74,73,72,72,73,74,76,76,76,76,76,76,76,76,76,76,76,76,76,74,73,72,72,72,70,68,65,64,62,61,60,60,60,60,60,58,58,58,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,61,62,64,64,62,62,62,64,64,64,64,64,64,64,64,64,64,64,64,64,62,61,60,58,57,56,57,58,60,60,60,60,58,57,56,56,54,53,50,49,48,49,52,54,56,56,56,56,56,56,56,56,56,56,56,56,56,54,52,50,50,50,49,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,49,50,52,52,52,50,49,49,50,50,49,48,48,48,46,45,44,44,44,44,44,44,44,44,42,42,42,44,44,44,44,44,44,44,44,44,44,44,44,44,44,44,44,44,44,44,44,42,41,40,40,40,40,40,38,37,36,36,34,33,32,32,32,33,34,36,36,36,36,34,33,32,32,32,32,32,32,32,32,32,32,32,32,33,34,36,36,36,36,36,36,37,38,40,41,42,44,44,45,46,49,50,52,52,52,52,52,52,50,49,48,48,48,48,48,48,48,48,48,48,46,45,44,44,42,41,40,40,40,40,41,42,44,44,44,44,44,44,44,45,46,49,50,52,52,52,52,52,52,52,53,54,56,56,56,56,56,56,56,56,56,56,56,56,56,57,60,62,64,64,64,64,64,64,64,64,64,64,62,61,60,58,57,56,56,56,56,56,56,54,54,56,58,61,62,64,62,61,60,60,60,60,60,60,60,60,60,60,60,60,61,62,65,66,68,68,68,68,69,70,72,72,72,72,72,72,72,72,72,72,70,69,68,68,66,65,64,64,64,64,62,61,60,60,60,60,60,60,60,60,60,58,57,56,56,56,56,56,57,57,57,54,52,49,48,48,49,50,52,52,52,52,52,52,52,52,52,50,49,48,46,45,44,44,45,46,46,46,46,48,48,48,48,48,49,50,52,52,52,52,52,52,52,50,49,48,48,48,48,48,48,48,48,49,50,52,52,52,52,52,50,49,48,48,48,48,48,48,48,49,50,52,52,52,52,52,52,52,52,52,52,52,52,50,49,48,46,45,44,42,41,40,38,36,33,32,32,32,32,32,32,32,32,32,32,33,34,36,34,33,32,30,29,26,25,24,24,24,22,22,22,24,24,25,26,28,26,25,24,24,22,21,20,20,20,20,20,20,21,22,24,24,24,24,24,22,22,22,24,24,24,22,21,20,20,20,20,20,20,20,20,20,20,20,20,18,17,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,14,13,12,10,9,8,8,6,5,4,5,6,8,6,5,4,4,4,4,4,4,4,5,8,12,14,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,17,18,20,20,20,20,20,18,17,16,16,16,16,16,14,12,9,8,8,8,8,6,5,4,4,4,4,4,4,4,4,4,4,5,5,5,4,4,5,5,5,4,5,5,5,4,3,3,3,4,4,4,4,4,4,4,4,4,4,4,5,5,5,3,3,4,5,6,8,8,9,10,12,12,12,12,12,12,12,10,9,8,8,8,8,8,8,6,6,5,5,4,5,6,8,8,8,8,8,8,8,8,8,8,6,5,4,4,4,4,5,6,8,8,8,6,5,4,4,4,5,6,8,8,9,10,12,12,10,10,12,14,14,13,12,12,12,12,12,12,12,12,12,12,12,12,10,9,8,8,8,8,8,8,8,8,9,10,12,12,13,14,16,16,16,14,13,12,13,16,18,20,21,22,22,21,20,20,20,20,20,20,20,20,20,20,18,18,18,20,20,20,20,20,20,18,17,16,16,16,16,16,14,13,12,12,12,12,12,12,12,10,9,8,8,8,8,9,10,12,10,9,8,8,8,9,10,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,14,16,16,16,14,13,12,12,12,12,12,10,10,10,10,9,8,8,9,9,9,6,5,4,4,4,4,4,4,4,4,4,4,4,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,6,9,10,13,14,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,17,18,20,20,20,20,20,20,20,18,17,17,18,20,20,20,20,20,20,20,20,20,18,17,14,12,9,8,8,9,10,12,13,14,16,14,14,14,16,14,13,12,10,9,8,8,6,5,4,4,5,6,8,8,6,5,4,4,4,4,4,4,4,3,3,3,4,4,4,4,4,5,8,9,9,6,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,3,3,3,4,3,3,3,4,4,5,5,5,4,5,6,8,6,5,5,6,8,8,8,8,8,8,8,8,8,6,5,4,4,4,4,4,5,7,7,7,6,6,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,6,8,8,6,5,5,6,8,9,10,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,14,16,16,16,17,18,20,20,20,20,20,20,20,20,18,18,18,20,20,20,18,17,16,16,16,16,16,16,16,16,14,13,12,13,14,17,18,20,18,17,14,13,12,12,12,12,12,12,12,12,10,9,8,8,8,8,6,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,7,6,8,6,5,4,4,4,4,4,4,4,4,4,4,5,8,10,13,14,16,16,16,17,18,20,20,20,20,21,22,24,24,22,21,20,20,20,18,17,16,16,16,16,14,13,12,13,14,16,16,16,16,16,16,16,16,16,17,18,20,20,20,21,22,24,24,24,25,26,28,28,28,29,30,32,32,32,30,29,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,26,25,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,22,21,20,20,20,20,18,17,16,16,16,16,14,13,12,13,14,14,13,12,10,9,8,8,8,9,10,12,12,12,12,12,10,8,7,5,5,4,5,8,10,12,12,12,12,12,12,13,14,16,16,16,16,17,18,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,21,22,24,24,25,25,25,24,24,24,24,24,25,26,26,24,21,20,20,20,20,21,22,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,22,21,20,20,20,20,21,22,24,24,24,24,22,21,20,20,21,22,24,24,24,24,25,25,25,24,22,21,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,18,17,16,16,16,16,16,16,16,16,16,17,18,20,20,18,17,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,17,18,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,18,17,14,14,14,16,16,16,16,16,14,14,14,16,16,16,16,16,16,16,16,16,14,13,12,12,12,13,14,17,18,20,20,20,18,17,16,16,14,13,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,12,12,12,10,9,8,8,8,8,8,8,8,8,8,8,8,8,9,12,13,14,14,16,16,16,14,12,9,8,8,8,6,5,4,4,5,6,8,8,8,8,8,8,8,8,8,8,8,8,8,9,10,12,12,12,12,13,14,16,16,14,13,12,12,12,12,13,14,16,16,16,16,16,16,16,16,17,18,20,20,20,20,20,20,20,18,17,16,16,16,14,13,12,12,12,12,12,10,8,5,4,4,4,4,4,4,4,4,3,2,1,2,3,4,3,4,6,8,8,8,8,8,8,8,8,8,8,8,6,6,8,10,12,12,12,12,12,12,12,13,13,13,12,12,12,12,12,10,9,6,6,4,6,6,8,8,8,6,5,4,4,3,4,4,5,4,4,4,4,4,4,5,5,5,4,4,4,5,8,10,10,9,8,8,6,5,4,4,4,5,5,5,5,6,8,8,8,8,8,8,8,8,8,8,8,8,6,5,4,4,4,4,5,6,8,8,6,5,4,4,4,4,5,6,8,8,8,8,8,9,10,12,12,12,12,12,12,10,9,8,9,12,14,16,16,17,18,18,17,16,16,17,18,20,20,20,20,20,20,20,20,20,20,18,17,16,16,16,16,16,16,16,16,16,16,16,16,17,18,18,17,16,16,14,13,12,12,12,12,12,12,12,10,10,9,9,8,8,8,8,8,9,10,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,9,8,8,8,8,8,8,8,6,5,4,4,5,5,7,7,8,8,8,9,10,12,12,12,12,12,12,12,12,12,12,12,13,14,17,18,20,18,17,16,16,17,17,18,18,20,20,20,21,21,21,18,18,18,20,20,18,17,16,16,16,16,16,14,13,13,14,14,13,12,12,12,12,12,10,9,8,8,8,8,8,8,8,6,5,4,4,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,4,4,5,6,8,8,8,8,9,10,12,12,13,14,16,17,18,18,17,16,16,16,14,13,12,12,12,12,12,12,12,12,12,12,10,9,8,8,8,8,6,6,6,8,8,9,10,12,13,16,18,20,20,18,17,16,16,16,16,16,16,16,14,13,12,12,12,10,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,5,5,5,5,4,3,3,3,4,5,7,8,6,5,4,4,4,5,6,6,7,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,6,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,10,12,12,12,10,9,8,8,8,8,8,8,8,8,8,9,10,12,12,12,12,12,12,13,16,18,20,20,20,18,17,16,16,16,16,17,18,20,20,20,18,17,16,14,13,12,12,12,12,13,13,13,13,14,16,16,16,16,16,16,16,16,16,14,13,12,12,12,10,9,9,9,9,8,8,8,8,8,6,6,4,4,4,4,4,3,5,6,8,8,8,8,8,6,5,5,5,5,4,4,4,4,4,4,4,4,5,6,8,8,8,8,8,8,8,8,8,9,10,12,12,12,12,12,12,12,12,12,10,9,8,6,5,5,6,8,8,9,10,13,16,18,20,20,20,21,21,21,20,20,20,21,22,24,25,26,28,28,28,29,30,32,32,32,32,32,33,34,36,36,36,36,36,36,36,36,36,36,34,32,29,28,28,28,28,28,28,28,26,25,24,24,24,24,24,24,24,24,22,21,18,17,16,16,16,16,16,16,16,16,16,16,16,16,17,18,20,20,20,20,20,20,20,20,18,17,17,18,21,22,24,24,24,24,24,22,21,20,20,20,20,20,20,20,20,18,17,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,14,13,10,9,6,5,4,4,4,4,4,4,4,4,4,4,5,6,8,8,8,6,5,4,5,5,5,4,4,5,6,8,8,8,8,8,6,5,4,5,6,6,5,5,5,5,4,4,4,4,4,4,4,4,4,4,5,8,10,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,9,8,6,5,4,5,6,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,5,4,4,4,4,5,6,8,8,8,8,8,8,8,8,8,6,5,5,6,9,10,10,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,10,10,12,12,12,12,12,12,12,12,12,12,10,9,8,8,8,8,8,9,10,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,14,16,16,16,16,16,16,14,13,12,13,14,16,16,16,16,16,16,16,16,17,18,20,20,20,20,20,20,20,20,20,20,18,17,17,18,20,20,18,16,13,12,12,12,12,12,12,12,12,12,12,12,13,13,13,12,12,12,12,12,12,13,14,16,16,16,16,16,14,13,13,14,16,14,13,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,12,12,12,12,12,13,14,16,16,14,13,12,10,10,9,9,8,8,8,8,8,8,8,8,9,10,12,12,12,12,12,12,12,12,13,14,17,18,20,20,20,20,20,20,20,20,18,17,14,13,12,12,12,12,12,10,9,6,5,4,4,4,4,4,4,4,4,3,3,3,4,4,5,6,8,8,6,5,4,4,5,6,8,8,8,8,6,5,4,4,4,4,4,4,4,4,4,5,6,8,8,8,8,8,9,10,12,12,12,12,12,12,10,9,8,8,8,8,9,10,12,13,14,17,18,20,20,20,20,20,20,20,18,17,16,16,14,13,10,9,8,8,8,8,8,8,8,9,10,12,12,10,9,8,8,8,8,6,5,4,4,4,4,3,3,3,4,4,4,4,6,7,8,8,8,8,8,8,8,8,8,6,5,4,4,4,5,6,8,9,10,10,9,8,8,8,8,6,5,4,4,5,6,6,4,3,3,4,4,4,4,4,4,5,5,5,4,5,6,6,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,6,8,8,8,8,9,10,12,12,12,12,12,12,12,12,10,9,8,8,8,8,8,8,9,10,12,12,12,12,13,14,16,17,18,18,17,17,18,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,21,22,24,24,24,24,25,26,28,29,30,32,32,32,32,32,32,33,34,36,34,32,29,28,28,28,28,29,30,32,32,33,34,36,36,34,34,36,40,41,41,40,40,40,40,40,40,38,36,33,32,32,32,30,30,30,32,32,32,32,32,32,32,32,32,30,29,28,28,28,26,25,24,24,24,24,22,21,18,16,13,13,14,16,16,17,18,20,20,20,20,20,20,21,22,24,24,24,24,24,24,24,22,21,20,20,20,18,18,18,18,16,13,12,12,12,12,12,12,12,12,12,12,10,9,8,8,9,9,9,8,8,8,9,10,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,14,16,18,20,20,21,22,24,24,24,24,24,24,24,24,24,24,25,26,28,28,28,28,28,28,28,28,28,28,29,30,32,32,30,29,28,29,30,32,30,29,29,30,30,29,28,28,28,29,32,36,40,42,44,44,44,44,44,44,44,44,45,48,50,52,52,52,52,52,52,52,52,50,49,48,48,48,46,45,44,44,44,45,46,48,48,48,48,48,48,48,48,48,46,44,41,40,40,40,40,40,40,41,42,44,44,44,42,41,40,40,40,40,40,38,37,36,36,36,36,36,37,38,40,40,40,40,40,40,40,40,40,41,42,44,44,44,45,46,48,48,48,48,48,49,49,49,48,48,48,48,48,48,48,48,48,48,48,48,48,49,50,52,52,52,50,49,48,48,48,48,48,48,48,48,48,48,48,49,50,52,52,52,52,52,52,52,52,52,50,49,46,45,45,46,48,48,48,46,46,46,48,48,48,49,50,52,52,52,52,52,52,52,52,52,53,54,56,56,54,53,52,52,52,53,54,56,56,56,56,56,56,56,56,57,58,60,60,60,60,60,60,60,60,58,57,56,56,56,56,56,56,57,58,60,60,60,60,60,60,61,64,66,68,68,68,66,65,62,61,60,58,57,56,56,56,56,56,56,56,56,56,56,56,56,54,53,52,52,52,50,49,48,48,48,48,48,48,48,48,48,48,48,48,48,48,49,50,52,52,52,52,52,52,52,52,52,52,52,52,52,52,52,53,54,56,56,56,57,58,60,60,60,60,60,60,60,61,61,61,60,60,60,60,60,60,60,61,62,64,64,64,64,65,65,64,60,56,53,52,52,53,54,56,56,56,56,56,56,56,54,53,52,52,52,52,52,52,53,54,56,56,56,56,56,56,57,58,60,60,60,60,58,58,57,56,54,54,56,56,56,56,56,56,56,56,56,56,56,56,57,58,60,60,60,60,60,60,60,60,60,60,60,60,60,60,61,62,64,64,64,64,64,64,64,64,62,61,60,60,58,57,56,56,56,56,56,56,57,58,60,61,62,64,64,64,64,64,64,64,64,64,64,65,66,69,70,72,72,70,69,66,65,64,64,64,64,62,62,62,64,64,64,64,62,61,60,60,60,60,60,60,60,60,60,58,57,56,56,54,53,52,53,53,53,52,52,52,52,52,53,54,56,54,53,52,52,52,52,52,53,54,56,54,53,52,52,52,52,52,52,52,50,49,48,46,45,44,44,44,44,44,44,44,42,41,41,42,44,45,46,48,48,48,48,48,48,48,48,48,49,52,54,56,56,56,57,58,60,60,60,60,60,60,60,60,60,60,60,60,60,60,58,57,56,56,56,57,58,60,61,62,64,64,64,62,61,60,60,60,60,60,61,62,64,64,64,64,64,65,66,68,68,68,68,68,68,69,70,72,72,72,73,74,76,76,76,76,74,73,72,72,72,72,72,70,70,70,70,68,65,65,65,65,62,60,57,56,56,56,56,56,56,54,53,52,52,52,52,52,52,52,50,50,50,52,52,53,54,56,57,60,62,62,61,60,60,60,58,57,56,56,56,56,56,56,56,56,54,53,52,52,52,52,50,49,48,48,48,48,46,45,44,44,44,44,44,44,44,44,44,45,45,45,44,44,44,44,44,44,42,41,40,40,40,41,42,44,44,44,44,45,46,48,48,48,49,50,50,50,50,52,52,52,53,54,56,54,54,54,56,56,56,56,56,56,56,56,56,56,56,54,53,52,52,53,54,56,56,56,56,56,56,56,57,58,60,60,61,62,64,64,64,64,64,65,66,68,68,69,70,72,72,72,72,72,72,72,72,72,72,72,72,72,72,72,72,72,72,72,72,72,70,69,68,68,68,68,68,68,68,68,68,68,68,68,68,68,66,65,64,64,64,64,64,62,62,62,65,66,68,66,65,64,64,62,61,60,60,60,60,60,60,60,60,60,60,60,60,60,61,62,64,64,64,65,65,65,64,64,64,64,64,64,64,62,62,62,64,62,62,62,64,64,64,64,64,64,62,61,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,61,61,61,60,60,60,60,60,60,60,61,62,64,65,66,68,68,69,70,72,72,72,72,72,72,72,72,72,72,72,72,72,72,72,72,72,70,68,65,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,62,61,60,60,60,60,60,60,58,57,56,56,56,56,56,56,56,56,54,52,50,50,52,52,52,53,54,56,56,54,52,49,48,48,48,48,48,46,46,46,48,49,50,52,52,52,52,52,52,52,53,54,54,53,52,52,52,52,52,52,52,52,52,52,52,52,53,54,56,56,56,57,57,57,56,56,56,56,56,56,54,53,52,53,54,56,56,56,56,54,53,52,52,52,52,52,50,49,48,48,48,46,45,44,44,45,46,48,48,48,48,48,48,48,48,48,48,48,48,46,45,45,46,48,48,48,46,45,44,44,44,45,46,48,48,48,49,50,53,53,53,52,50,49,46,45,42,41,40,40,40,40,38,36,33,32,32,32,32,32,33,34,34,32,29,28,28,28,28,29,30,32,32,32,32,32,32,32,32,32,32,33,34,36,36,36,34,33,32,32,33,34,36,36,36,36,37,37,38,38,40,40,40,40,40,40,41,42,44,44,44,44,44,42,41,40,40,40,38,37,36,36,36,36,36,36,36,36,36,36,37,38,40,40,40,41,42,42,41,40,40,40,40,40,40,40,41,41,41,40,40,40,40,40,40,38,37,36,36,36,36,36,36,36,37,38,41,42,44,44,44,45,46,46,45,44,44,44,44,44,44,44,44,45,46,48,48,48,48,48,48,48,48,49,50,52,52,53,54,56,56,56,54,52,49,48,48,48,48,48,48,48,48,46,45,44,44,44,44,44,44,44,44,44,44,44,45,46,48,46,45,44,44,45,48,50,52,50,48,45,44,44,44,44,44,44,44,42,41,40,40,40,40,40,40,40,40,40,40,40,40,40,40,40,38,37,36,34,33,33,34,34,32,29,28,29,30,32,32,32,32,32,33,34,36,36,36,36,36,36,36,34,32,28,25,25,25,25,24,24,24,22,20,17,16,17,18,20,20,20,20,21,22,24,24,22,21,20,18,17,16,16,16,16,14,13,12,12,13,14,16,17,18,20,20,20,20,20,20,20,20,20,20,18,17,16,16,16,17,18,20,20,20,20,20,20,20,20,20,20,20,20,20,18,17,16,16,16,16,16,16,16,16,14,13,12,10,9,8,8,8,8,8,8,9,10,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,14,16,16,16,16,16,16,16,16,14,13,12,12,12,12,12,12,12,12,10,9,8,8,6,5,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,4,4,4,4,4,5,6,8,6,5,4,4,4,4,4,4,4,4,4,4,4,4,4,5,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,6,8,8,8,8,8,8,9,9,9,8,8,8,8,8,8,9,10,12,10,9,8,8,8,8,8,8,8,8,9,10,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,16,18,20,21,22,24,24,24,24,25,26,26,25,24,24,22,21,20,20,18,17,16,16,16,16,16,16,16,16,17,18,20,20,20,20,20,20,20,18,17,17,18,20,20,20,20,20,20,20,20,21,21,20,17,16,16,16,16,16,17,17,17,16,16,16,16,16,16,16,16,16,16,14,13,12,13,14,16,16,16,16,14,13,12,12,12,12,12,12,12,10,9,8,8,8,8,8,8,8,8,6,5,4,4,4,4,4,4,4,4,4,4,4,4,4,5,6,6,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,6,8,6,6,5,5,4,4,4,4,4,4,4,4,3,3,4,5,5,4,4,4,4,5,8,10,12,10,9,8,8,8,8,9,10,12,12,12,10,9,6,5,5,6,8,8,8,8,8,8,8,8,8,8,8,8,8,6,5,4,4,4,4,5,6,8,8,8,6,5,4,4,4,4,4,4,4,4,5,6,8,8,8,8,8,8,6,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,6,8,8,9,10,12,12,12,12,13,14,17,18,20,20,20,20,21,22,24,24,24,24,24,24,24,22,21,20,20,20,20,20,20,20,20,20,20,20,18,17,16,16,16,16,16,16,16,16,16,17,20,22,24,25,26,28,28,28,28,28,28,28,29,30,32,32,30,30,30,32,32,32,32,32,32,32,32,30,29,26,25,24,24,24,22,21,20,20,20,20,20,20,20,18,17,16,16,16,17,18,20,20,20,20,20,20,20,20,20,20,21,22,22,21,20,20,18,17,16,16,14,13,12,12,13,14,16,16,16,16,16,16,16,16,14,13,12,12,10,9,8,8,8,8,8,6,5,4,4,4,5,6,8,9,10,12,10,9,9,9,9,8,6,5,4,4,4,4,5,6,8,6,5,4,4,6,8,10,12,12,12,12,12,13,14,16,16,16,16,16,16,16,16,16,16,16,16,16,16,14,13,12,12,12,12,12,10,9,8,8,8,8,8,8,8,8,8,8,6,5,4,4,5,5,5,4,5,5,5,4,4,4,4,5,6,8,8,8,8,6,5,4,4,4,4,5,6,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,10,10,9,8,8,8,8,8,8,9,10,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,12,12,12,12,13,14,16,16,16,16,16,17,18,18,17,16,16,16,14,13,12,12,13,14,16,16,16,16,16,16,16,16,16,14,13,12,12,12,12,13,14,16,16,16,16,16,16,16,17,18,18,17,16,16,16,16,16,16,16,16,16,17,18,20,18,17,16,16,14,13,12,12,12,13,14,16,16,16,17,18,20,20,20,18,18,18,18,18,18,20,20,21,22,24,24,22,20,17,16,16,16,16,14,13,12,12,12,12,12,12,12,12,13,14,16,16,16,16,16,16,16,16,16,16,16,16,16,17,17,17,16,17,18,20,18,17,16,16,16,14,13,12,12,12,12,12,12,10,9,8,8,8,8,8,9,10,12,12,12,12,12,12,12,10,9,8,9,10,12,12,12,10,9,8,8,8,8,8,8,8,8,8,8,8,8,8,6,5,4,4,5,6,8,8,8,6,5,4,5,8,10,13,14,14,13,12,12,12,12,12,13,14,16,16,16,16,16,14,14,14,14,13,12,12,12,12,10,8,5,4,4,3,4,5,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,5,4,5,6,9,12,13,13,12,10,9,8,8,8,8,6,5,5,6,8,8,8,8,8,6,5,4,4,4,4,4,4,3,3,3,3,5,5,6,6,8,8,8,8,8,6,5,4,4,4,4,4,5,6,8,8,6,5,4,4,4,4,4,4,4,3,3,3,4,3,4,4,3,3,2,3,3,4,5,8,10,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,14,16,16,14,13,12,13,16,18,20,21,22,24,24,24,22,21,20,21,22,24,22,21,20,20,20,18,17,16,16,16,16,16,16,16,16,16,16,16,16,16,14,13,12,13,14,16,14,14,14,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,14,12,9,8,8,8,8,8,8,8,8,8,8,8,8,9,10,12,12,12,12,12,12,12,12,12,12,12,12,12,13,14,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,14,13,12,12,12,12,12,12,13,13,12,9,8,8,8,8,8,8,8,8,8,8,8,9,10,13,14,14,13,12,12,12,10,9,9,10,12,12,12,13,14,14,13,12,12,12,12,12,12,12,13,16,18,20,20,20,20,18,17,16,16,16,16,16,16,16,17,18,20,20,20,20,20,20,20,20,20,20,20,20,20,20,18,16,13,12,12,12,10,9,9,12,14,16,17,18,20,20,20,20,20,20,20,21,22,22,21,20,20,18,17,16,17,18,20,20,21,22,24,24,24,24,24,24,24,24,25,26,28,28,28,28,28,28,28,28,29,30,32,32,32,32,32,32,30,29,28,28,28,28,28,29,30,32,32,32,33,34,37,40,42,44,44,44,42,41,40,40,40,40,40,40,40,40,40,40,40,40,40,40,40,40,40,40,40,40,40,40,40,40,40,41,42,44,44,44,44,44,44,42,41,40,40,38,37,36,36,36,36,36,36,36,36,34,34,34,34,33,32,32,32,32,32,32,32,30,29,28,26,25,24,24,24,24,24,24,24,22,21,20,20,18,17,16,16,16,17,18,20,20,20,21,22,24,24,24,25,26,26,25,24,24,22,21,20,20,20,20,20,18,17,16,16,16,16,16,16,17,17,17,16,16,16,16,16,16,16,16,16,14,13,10,9,6,5,4,5,6,8,8,9,10,12,12,12,12,12,13,14,16,16,17,18,20,20,18,17,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,17,18,20,21,22,24,24,24,24,24,22,21,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,21,22,25,26,28,28,29,30,32,33,36,38,40,40,40,40,40,40,40,40,41,42,44,44,44,44,44,44,44,44,44,44,45,46,48,48,46,45,44,45,46,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,49,50,52,52,53,54,56,56,56,56,56,56,56,56,56,56,56,56,56,56,57,58,61,62,64,62,62,61,61,60,60,60,60,60,58,57,57,58,60,60,60,60,60,60,60,61,62,64,64,64,64,64,64,64,64,64,64,64,65,65,65,62,61,60,60,58,56,53,53,54,56,56,56,56,56,56,56,56,57,58,60,60,60,60,60,60,60,60,60,60,58,57,56,54,52,49,48,48,48,48,49,50,53,54,54,53,52,52,53,53,54,54,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,54,54,53,53,53,54,56,56,56,56,57,58,60,60,60,60,60,60,60,60,60,60,60,58,57,56,54,52,50,50,52,52,52,52,53,54,56,56,56,56,56,56,57,60,62,62,61,60,60,60,58,57,56,56,56,56,57,57,56,53,52,52,52,53,54,54,54,54,56,56,56,56,56,56,57,58,60,60,58,57,56,56,56,56,56,56,56,56,56,57,57,57,56,56,54,53,52,52,52,52,52,52,52,52,52,52,52,52,52,50,49,48,48,48,48,48,46,45,44,45,46,49,50,52,52,50,49,49,52,54,56,57,58,60,60,60,60,60,60,58,57,56,56,56,56,56,56,56,56,56,56,54,53,52,52,53,54,56,56,56,56,56,56,57,60,64,66,68,68,68,68,68,68,68,66,65,65,66,68,68,68,68,68,68,68,68,68,68,68,66,65,64,64,64,65,66,68,68,66,65,64,64,62,61,60,60,60,60,60,58,57,56,54,54,54,56,56,56,56,56,56,56,56,57,60,62,64,64,64,64,64,64,64,64,64,64,65,66,68,68,68,68,68,68,68,68,66,64,61,60,60,60,60,61,62,64,64,64,65,66,68,68,68,68,68,68,69,70,73,74,76,76,76,77,78,80,80,80,80,80,80,78,77,76,76,76,76,76,76,76,76,76,74,73,72,72,70,69,69,70,72,72,72,72,72,72,72,72,72,73,74,76,76,76,76,77,78,80,81,82,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,85,86,89,90,92,92,92,90,88,85,84,82,81,81,82,84,84,84,84,84,84,84,84,84,84,84,84,84,82,81,78,77,76,77,77,77,76,76,77,80,81,81,80,80,80,80,80,80,80,80,80,80,78,77,76,76,77,78,80,80,81,84,86,88,88,88,88,88,88,86,85,84,84,84,84,84,84,84,84,84,82,81,80,80,80,81,84,86,88,88,88,88,89,90,92,92,92,92,92,92,93,94,94,93,92,92,92,92,93,94,96,96,96,96,96,96,96,96,96,96,96,96,96,96,94,94,94,96,96,96,96,97,98,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,98,97,96,96,96,97,98,100,100,100,100,100,100,100,100,100,100,100,100,100,100,98,97,96,94,93,92,92,92,92,92,92,92,92,92,92,92,92,92,92,92,90,89,86,85,84,84,84,84,82,81,80,80,81,82,84,84,84,82,81,80,80,80,80,80,80,80,80,80,80,80,80,80,81,81,82,81,80,77,76,76,74,73,70,69,68,68,69,70,72,70,69,68,68,68,68,68,68,68,68,68,69,72,74,76,76,74,72,69,69,69,69,68,68,68,66,65,65,66,68,68,68,68,68,69,70,72,72,72,72,72,72,72,73,74,76,76,76,76,76,76,76,76,76,76,76,74,73,72,72,73,74,76,76,77,78,80,80,80,80,80,80,80,80,78,77,76,76,76,74,73,72,72,73,74,76,76,76,76,76,76,76,76,76,76,76,76,76,76,76,76,77,78,80,80,80,80,80,78,77,74,73,72,72,72,73,76,78,80,78,78,78,80,80,80,80,80,78,77,76,74,73,72,72,72,72,72,72,72,70,69,68,68,68,68,68,66,64,61,61,64,68,70,70,69,68,68,68,69,70,72,72,72,70,69,68,68,68,68,69,70,72,72,72,72,72,72,72,72,70,69,68,68,68,68,68,68,68,68,66,65,64,64,64,64,64,64,64,64,64,64,62,61,60,60,58,57,56,57,58,60,60,60,60,60,60,60,60,60,60,60,61,62,64,62,61,60,60,60,60,60,58,57,56,54,53,52,52,52,52,52,52,52,52,52,52,52,52,52,52,53,54,57,58,60,60,60,60,60,60,60,60,60,58,57,56,56,56,57,57,57,56,56,56,56,57,58,58,57,56,56,57,58,60,60,58,57,56,56,56,56,56,56,54,53,52,52,52,52,52,52,52,52,52,53,54,56,56,54,53,52,52,52,50,49,48,48,48,48,48,48,46,44,42,41,41,40,40,41,42,44,44,44,44,42,41,40,40,40,40,40,40,40,40,41,42,44,44,44,44,45,46,48,48,48,48,49,50,52,53,54,56,56,56,57,58,60,61,62,65,66,68,66,65,64,64,64,64,64,64,64,64,65,66,68,68,68,68,68,69,69,69,69,70,72,72,72,72,70,69,68,68,68,68,68,68,68,68,69,70,72,72,72,72,72,72,72,72,72,72,72,73,74,76,74,73,70,69,68,68,68,68,68,68,68,68,68,68,68,66,66,66,68,68,69,70,72,72,72,72,72,70,69,68,68,68,68,68,69,70,72,72,72,72,72,72,70,69,68,69,69,70,70,70,69,68,68,68,68,68,68,66,65,64,64,64,65,66,68,68,68,68,68,66,66,66,68,68,68,68,68,68,68,66,65,64,64,64,62,61,60,60,60,58,57,56,54,53,52,52,50,49,46,45,45,46,48,48,48,46,45,44,45,46,48,46,45,44,44,44,44,44,44,44,44,44,44,44,44,44,44,44,44,42,41,40,40,40,40,40,40,40,41,42,45,46,48,48,48,48,48,48,48,48,48,48,48,48,48,48,46,45,44,44,42,41,40,38,37,36,36,36,36,36,36,36,36,36,36,36,36,36,36,34,34,34,36,34,33,32,30,29,29,30,32,32,32,32,32,30,29,28,28,28,28,28,26,24,21,20,18,17,17,18,20,18,17,16,16,16,16,14,13,12,12,10,10,10,10,9,8,8,8,8,8,8,8,8,8,8,6,5,4,4,4,4,4,4,5,5,5,4,4,4,4,4,4,4,4,4,4,3,3,3,4,4,4,4,4,4,4,4,4,4,4,5,6,8,8,6,5,4,4,4,4,4,4,4,4,4,4,4,6,7,9,10,12,12,12,12,12,12,12,12,12,13,14,16,16,16,16,16,16,16,14,13,12,12,12,12,13,14,16,16,16,16,16,16,16,17,18,20,20,20,20,20,20,20,20,20,20,20,20,20,18,17,17,18,20,20,20,20,20,21,22,24,24,24,24,24,24,22,20,17,16,16,16,14,12,9,8,8,8,8,8,8,8,8,9,10,12,12,12,13,14,16,16,16,16,16,17,18,20,20,20,20,18,17,16,16,17,18,20,20,20,20,20,20,20,20,20,20,20,20,20,20,21,22,24,24,24,24,24,24,24,22,21,20,20,20,20,20,20,18,17,14,13,12,12,13,14,16,16,16,14,14,14,16,16,16,16,16,16,16,16,16,17,18,20,20,20,20,20,20,20,21,22,24,24,24,24,24,24,24,24,24,22,21,20,20,20,20,20,20,18,17,16,16,16,16,16,16,16,16,16,17,18,20,20,20,20,20,20,20,20,20,20,20,20,20,20,21,22,24,24,24,24,24,24,25,26,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,26,25,24,25,26,28,28,28,28,28,28,28,29,30,32,32,32,32,32,32,32,32,32,32,32,32,32,32,32,32,32,32,32,32,32,32,30,29,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,26,25,24,24,24,25,28,30,32,30,29,28,28,28,28,28,28,28,29,29,29,28,28,28,28,29,30,32,32,32,32,33,34,36,37,38,40,40,40,40,41,42,44,44,44,44,44,45,46,48,48,46,45,44,44,44,44,42,42,42,44,44,44,44,42,41,41,42,44,45,46,48,48,48,49,50,52,50,49,46,45,44,44,44,44,44,44,42,41,40,40,40,40,40,40,40,40,40,40,40,40,41,42,44,44,44,44,44,44,44,44,44,44,44,42,41,40,40,40,40,40,40,40,40,38,37,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,34,33,32,32,32,32,32,32,32,32,30,28,25,24,24,25,28,30,32,32,32,32,32,32,32,33,33,33,32,32,32,30,29,28,28,28,28,29,29,29,28,28,28,26,25,24,24,24,24,24,24,22,21,20,21,22,24,24,24,24,25,28,30,32,32,32,33,36,38,41,42,44,42,41,40,41,42,45,46,48,48,48,48,48,46,45,44,44,44,44,42,41,40,40,40,40,40,40,40,40,40,40,40,40,40,40,40,40,38,37,36,36,36,36,36,36,36,36,36,37,40,42,44,44,44,44,44,44,44,44,44,42,41,41,42,44,44,44,44,44,44,44,44,44,44,44,45,46,49,50,52,52,50,50,50,52,52,50,49,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,49,50,52,52,53,54,54,53,53,54,56,56,56,56,56,57,58,60,60,60,60,60,61,64,66,69,72,74,76,76,76,76,76,76,76,76,76,76,76,76,76,77,78,80,80,80,80,80,80,81,82,82,81,80,80,80,80,80,78,77,77,78,80,80,80,80,80,78,77,76,77,78,80,80,80,80,78,78,78,80,80,80,80,80,80,81,84,86,88,88,88,88,88,88,88,86,85,85,86,86,86,86,88,86,85,84,84,84,85,86,88,88,88,86,85,84,85,86,88,88,88,88,88,88,86,85,84,84,84,84,85,86,86,85,84,84,84,85,86,86,84,81,80,81,82,84,84,84,84,84,84,84,82,81,81,82,84,82,81,78,77,76,76,76,77,78,80,80,81,82,84,84,84,84,82,82,82,82,81,80,80,80,78,77,76,74,73,72,72,73,74,76,77,78,80,80,80,80,80,80,80,80,78,77,76,76,76,76,77,78,80,80,80,80,80,81,82,84,84,84,84,84,84,84,84,84,84,84,84,84,84,82,81,80,80,80,80,80,80,80,81,82,85,88,90,92,92,93,94,96,96,96,96,97,98,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,98,97,96,96,96,96,96,94,93,92,92,90,89,88,88,89,90,92,92,93,96,98,100,100,100,100,100,100,98,98,98,100,100,100,98,96,93,92,92,92,92,93,96,98,100,98,97,96,96,97,98,100,100,100,98,96,93,92,92,92,90,89,88,88,88,88,88,88,86,85,84,84,82,81,80,80,80,80,80,80,81,82,84,84,84,85,86,88,88,88,88,89,90,92,92,92,92,90,89,88,88,88,88,88,88,88,88,88,88,86,85,84,85,86,88,88,88,88,88,88,88,88,88,88,88,88,88,88,88,88,88,88,88,88,88,88,86,85,85,86,86,85,84,84,82,81,80,80,80,80,80,80,80,80,78,78,78,80,80,80,80,80,80,80,80,80,80,80,78,77,76,76,74,73,72,72,72,73,74,76,77,78,80,80,80,80,80,80,80,80,80,81,81,81,80,78,77,76,76,76,76,76,76,76,76);




variable  height:  integer := 0 ;
variable index:  integer := 0 ;
variable counter : integer:= 0;
constant MaxNum : integer := 750000;
constant gap : integer := 360;
   

begin
	if RESETn = '0' then
	   mVGA_R <= "000" ;	
      mVGA_G <= "000" ;	
    mVGA_B <= "00" ;
		
		
		drawing_request	<=  '0' ;

		elsif rising_edge(CLK) then
		
		
		    if (index = 14722) then
			        index:=0;
		    end if;	
		
			if (counter=MaxNum) then
			     counter:=0;
			     index:=index+2; -- controlling speed
				  
			else 
			     counter :=counter +1;
			end if;
			
			

			 
			 	
			if (counter<MaxNum) then
			
			     height := height_value( index + oCoord_X); -- oCoord_X for 640 offset
				 
			   if (oCoord_Y < height+20 or  oCoord_Y>height+gap+20) then 
			
			   			mVGA_R <= "101" ;	
			            mVGA_G <= "101" ;	
			            mVGA_B <= "10" ;
							
						
			        drawing_request	<= '1'; 
				 else
							mVGA_R <= "000" ;	
			            mVGA_G <= "000" ;	
			            mVGA_B <= "00" ;
						
			        drawing_request	<= '0'; 
			    end if;
				 
				 
				
				
			end if;
			
			
			
			
	 
	end if;

  end process;

	
end behav;		