library IEEE;
use IEEE.STD_LOGIC_1164.all;
--use IEEE.std_logic_unsigned.all;
--use ieee.numeric_std.all;
--use ieee.std_logic_arith.all;
-- Alex Grinshpun April 2017
-- Dudy Nov 13 2017


entity obstacle_draw is
port 	(
		--////////////////////	Clock Input	 	////////////////////	
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		ObjectStartX	: in integer;
		ObjectStartY 	: in integer;
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0)

		
	); 
end obstacle_draw;

architecture behav of obstacle_draw is 

constant object_X_size : integer := 38;
constant object_Y_size : integer := 61;

--constant object_X_size : integer := 85;
--constant object_Y_size : integer := 30;



type ram_array_obstacle is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);  
  
constant object_colors_obstacle: ram_array_obstacle := ( 


(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"92",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"24",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"b6",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"b6",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"24",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"6d",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"24",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"b6",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"b6",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"24",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"49",x"24",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"24",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"6d",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"24",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"24",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"24",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"6d",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"24",x"6d",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"24",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"b6",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"b6",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"24",x"6d",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"24",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"6d",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"6d",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"24",x"6d",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"24",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"b6",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"b6",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"24",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"24",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"6d",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"24",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"24",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"24",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"6d",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"24",x"24",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"b6",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"b6",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"24",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"b6",x"6d",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"24",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"b6",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"b6",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"92",x"6d",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"24",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"24",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"24",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"24",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"24",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"24",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"b6",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"b6",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"6d",x"b6",x"b6",x"b6",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"24",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"24",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"6d",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"00",x"00",x"00",x"00",x"00")




);





-- one bit mask  0 - off 1 dispaly 
type object_form_obstacle is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object_obstacle : object_form_obstacle := (

("00000000000000000000000000000000000000"),
("00000000000000000000000000000000000000"),
("00000000000000000000000000000000000000"),
("00001111111111111111111111111111000000"),
("00001111111111111111111111111111100000"),
("00001111111111111111111111111111000000"),
("00001111111111111111111111111111000000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00001111111111111111111111111111100000"),
("00001111111111111111111111111111000000"),
("00001111111111111111111111111111000000"),
("00011111111111111111111111111111110000"),
("00111111111111111111111111111111110000"),
("00111111111111111111111111111111110000"),
("00111111111111111111111111111111110000"),
("00111111111111111111111111111111110000"),
("00011111111111111111111111111111100000"),
("00001111111111111111111111111111000000"),
("00001111111111111111111111111111000000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00001111111111111111111111111111000000"),
("00001111111111111111111111111111000000"),
("00001111111111111111111111111111100000"),
("00111111111111111111111111111111110000"),
("00111111111111111111111111111111110000"),
("00111111111111111111111111111111110000"),
("00111111111111111111111111111111110000"),
("00111111111111111111111111111111110000"),
("00001111111111111111111111111111000000"),
("00001111111111111111111111111111000000"),
("00001111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00001111111111111111111111111111000000"),
("00001111111111111111111111111111000000"),
("00001111111111111111111111111111100000"),
("00111111111111111111111111111111110000"),
("00111111111111111111111111111111110000"),
("00111111111111111111111111111111110000"),
("00111111111111111111111111111111110000"),
("00111111111111111111111111111111110000"),
("00001111111111111111111111111111000000"),
("00001111111111111111111111111111000000"),
("00001111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000"),
("00011111111111111111111111111111100000")



);





signal bCoord_X : integer := 0;-- offset from start position 
signal bCoord_Y : integer := 0;



signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';

--		
signal objectEndX : integer;
signal objectEndY : integer;


begin

-- Calculate object end boundaries
objectEndX	<= object_X_size+ObjectStartX;
objectEndY	<= object_Y_size+ObjectStartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

-- test if ooCoord is in the rectangle defined by Start and End 
	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectEndX) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectEndY) else '0';

-- calculate offset from start corner 
	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
 


process ( RESETn, CLK)



  	variable counter : integer:= 0;
   constant MaxNum2 : integer := 45000000;
	
	--- i want to print a picture every 750000
 	
   begin
	
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;

		
		elsif rising_edge(CLK) then
	
				mVGA_RGB	<=  object_colors_obstacle(bCoord_Y , bCoord_X);	
			   drawing_request	<= object_obstacle(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; 		

			
	end if;

  end process;

		
end behav;		
		