library IEEE;
use IEEE.STD_LOGIC_1164.all;
--use IEEE.std_logic_unsigned.all;
--use ieee.numeric_std.all;
--use ieee.std_logic_arith.all;
-- Alex Grinshpun April 2017
-- Dudy Nov 13 2017


entity cieling_object is
port 	(
		--////////////////////	Clock Input	 	////////////////////	
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		ObjectStartX	: in integer;
		ObjectStartY 	: in integer;
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0);
		MaxNum		: in integer
		
	);
end cieling_object;

architecture behav of cieling_object is 

constant object_X_size : integer := 640;
constant object_Y_size : integer := 200;
--constant R_high		: integer := 7;
--constant R_low		: integer := 5;
--constant G_high		: integer := 4;
--constant G_low		: integer := 2;
--constant B_high		: integer := 1;
--constant B_low		: integer := 0;





type ram_array1 is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);  

-- 8 bit - color definition : "RRRGGGBB"  
constant object_colors: ram_array1 := ( 


(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"04",x"04",x"00",x"08",x"08",x"00",x"04",x"08",x"04",x"04",x"35",x"35",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"08",x"35",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"08",x"35",x"2c",x"00",x"04",x"04",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"04",x"51",x"55",x"4d",x"28",x"55",x"55",x"24",x"2d",x"55",x"51",x"04",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"04",x"08",x"04",x"00",x"04",x"08",x"04",x"00",x"04",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"04",x"00",x"04",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"04",x"04",x"00",x"04",x"04",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"04",x"04",x"00",x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"04",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"04",x"00",x"04",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"00",x"00",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"00",x"00",x"04",x"08",x"00",x"00",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"4d",x"55",x"4d",x"00",x"00",x"00",x"00",x"00",x"24",x"55",x"55",x"04",x"08",x"35",x"35",x"35",x"00",x"04",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"04",x"00",x"00",x"08",x"08",x"04",x"00",x"04",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"51",x"55",x"04",x"08",x"35",x"2c",x"00",x"51",x"51",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"00",x"08",x"04",x"04",x"55",x"35",x"2d",x"28",x"55",x"55",x"24",x"2d",x"55",x"51",x"04",x"35",x"35",x"30",x"00",x"04",x"08",x"04",x"00",x"04",x"08",x"04",x"00",x"04",x"08",x"04",x"00",x"00",x"08",x"00",x"04",x"08",x"04",x"00",x"00"),
(x"00",x"00",x"00",x"2d",x"55",x"51",x"00",x"51",x"55",x"4d",x"00",x"4d",x"55",x"29",x"00",x"04",x"08",x"00",x"00",x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"55",x"24",x"00",x"08",x"04",x"00",x"00",x"00",x"00",x"4d",x"55",x"51",x"00",x"4d",x"75",x"4d",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"04",x"00",x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"00",x"00",x"08",x"08",x"00",x"04",x"08",x"04",x"00",x"00",x"00",x"00",x"04",x"08",x"04",x"00",x"08",x"04",x"00",x"29",x"55",x"04",x"00",x"00",x"00",x"00",x"51",x"4d",x"00",x"04",x"04",x"00",x"51",x"4d",x"00",x"4d",x"51",x"00",x"08",x"04",x"00",x"08",x"00",x"00",x"51",x"04",x"28",x"4d",x"00",x"04",x"00",x"04",x"04",x"00",x"04",x"00",x"2d",x"2d",x"00",x"00",x"00",x"04",x"08",x"00",x"04",x"71",x"24",x"00",x"08",x"00",x"28",x"75",x"24",x"00",x"08",x"04",x"00",x"08",x"00",x"00",x"28",x"00",x"2d",x"55",x"04",x"00",x"08",x"04",x"00",x"08",x"00",x"00",x"08",x"00",x"2d",x"51",x"00",x"00",x"00",x"00",x"04",x"00",x"04",x"00",x"04",x"71",x"00",x"28",x"51",x"00",x"2d",x"51",x"00",x"4d",x"51",x"00",x"00",x"00",x"00",x"00",x"08",x"04",x"00",x"4d",x"51",x"00",x"29",x"51",x"00",x"28",x"75",x"24",x"00",x"08",x"04",x"00",x"00",x"00",x"00",x"2d",x"51",x"00",x"4d",x"51",x"00",x"04",x"08",x"00",x"04",x"08",x"00",x"2d",x"51",x"00",x"04",x"08",x"00",x"00",x"00",x"00",x"04",x"08",x"00",x"04",x"08",x"00",x"00",x"00",x"00",x"04",x"04",x"04",x"51",x"00",x"4d",x"04",x"00",x"04",x"00",x"51",x"28",x"00",x"04",x"00",x"00",x"00",x"00",x"04",x"00",x"28",x"4d",x"00",x"4d",x"00",x"51",x"04",x"51",x"29",x"00",x"08",x"04",x"00",x"08",x"00",x"28",x"75",x"04",x"28",x"55",x"28",x"00",x"08",x"04",x"00",x"00",x"00",x"00",x"4d",x"51",x"00",x"4d",x"51",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"04",x"04",x"04",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4d",x"55",x"28",x"00",x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"04",x"04",x"08",x"08",x"00",x"04",x"08",x"08",x"04",x"04",x"55",x"55",x"28",x"00",x"51",x"55",x"28",x"04",x"55",x"51",x"00",x"04",x"08",x"00",x"24",x"55",x"55",x"04",x"00",x"08",x"08",x"04",x"00",x"08",x"08",x"00",x"28",x"75",x"28",x"00",x"08",x"04",x"00",x"29",x"75",x"51",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"4d",x"75",x"2d",x"00",x"04",x"08",x"04",x"28",x"75",x"29",x"00",x"08",x"08",x"00",x"28",x"55",x"51",x"00",x"00",x"08",x"08",x"04",x"00",x"08",x"08",x"04",x"00",x"00",x"00",x"00",x"04",x"55",x"4d",x"00",x"00",x"00",x"2d",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"04",x"55",x"55",x"04",x"08",x"35",x"35",x"35",x"00",x"28",x"55",x"51",x"00",x"04",x"08",x"08",x"04",x"00",x"51",x"55",x"51",x"00",x"28",x"55",x"55",x"4d",x"00",x"4d",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"00",x"4d",x"4d",x"00",x"04",x"08",x"00",x"04",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"00",x"28",x"51",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"08",x"04",x"04",x"08",x"08",x"00",x"04",x"08",x"08",x"00",x"04",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"51",x"75",x"28",x"00",x"00",x"00",x"00",x"31",x"55",x"04",x"08",x"35",x"2c",x"00",x"51",x"55",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"0c",x"24",x"55",x"51",x"04",x"35",x"35",x"2d",x"28",x"55",x"35",x"04",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"51",x"55",x"4d",x"28",x"55",x"55",x"4d",x"00",x"4d",x"55",x"51",x"00",x"24",x"75",x"04",x"28",x"75",x"2d",x"00",x"08"),
(x"28",x"28",x"00",x"2d",x"35",x"51",x"04",x"31",x"55",x"2d",x"00",x"2d",x"55",x"28",x"00",x"51",x"55",x"04",x"04",x"55",x"55",x"04",x"04",x"28",x"08",x"00",x"04",x"28",x"04",x"00",x"51",x"55",x"04",x"00",x"55",x"4d",x"00",x"08",x"28",x"00",x"2d",x"55",x"51",x"00",x"2c",x"55",x"2d",x"00",x"28",x"28",x"04",x"00",x"51",x"55",x"2d",x"00",x"08",x"28",x"28",x"00",x"04",x"28",x"28",x"00",x"4d",x"55",x"51",x"00",x"51",x"51",x"00",x"04",x"2c",x"04",x"04",x"55",x"55",x"04",x"04",x"55",x"51",x"00",x"28",x"55",x"51",x"00",x"28",x"28",x"00",x"28",x"55",x"28",x"00",x"55",x"51",x"00",x"2d",x"55",x"04",x"00",x"28",x"04",x"00",x"51",x"2d",x"00",x"4d",x"51",x"00",x"31",x"2d",x"00",x"2d",x"31",x"00",x"51",x"4d",x"04",x"55",x"24",x"00",x"51",x"04",x"28",x"2d",x"00",x"51",x"24",x"28",x"29",x"00",x"4d",x"00",x"2d",x"2d",x"00",x"28",x"00",x"28",x"55",x"04",x"04",x"55",x"04",x"28",x"55",x"04",x"28",x"55",x"04",x"04",x"55",x"2d",x"00",x"51",x"04",x"04",x"75",x"04",x"2d",x"55",x"04",x"24",x"55",x"28",x"24",x"55",x"24",x"04",x"51",x"00",x"2d",x"51",x"00",x"28",x"04",x"00",x"4d",x"00",x"4d",x"24",x"04",x"51",x"00",x"28",x"51",x"00",x"28",x"51",x"00",x"31",x"51",x"00",x"04",x"28",x"04",x"00",x"51",x"51",x"00",x"2d",x"51",x"00",x"2c",x"31",x"00",x"28",x"55",x"04",x"04",x"55",x"28",x"00",x"28",x"08",x"00",x"2d",x"31",x"00",x"2d",x"31",x"00",x"4d",x"51",x"00",x"4d",x"51",x"00",x"2d",x"55",x"00",x"29",x"55",x"00",x"00",x"28",x"00",x"28",x"55",x"04",x"28",x"51",x"00",x"04",x"04",x"00",x"51",x"28",x"00",x"51",x"00",x"4d",x"04",x"04",x"51",x"00",x"51",x"28",x"00",x"51",x"00",x"04",x"04",x"00",x"51",x"04",x"28",x"2d",x"00",x"4d",x"04",x"51",x"04",x"31",x"2c",x"00",x"51",x"28",x"00",x"51",x"04",x"28",x"55",x"04",x"28",x"55",x"28",x"00",x"51",x"2d",x"00",x"28",x"08",x"00",x"2d",x"51",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"24",x"55",x"55",x"04",x"2d",x"55",x"51",x"00",x"28",x"55",x"51",x"00",x"04",x"28",x"04",x"00",x"08",x"28",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4d",x"55",x"2d",x"00",x"08",x"28",x"00",x"00",x"00",x"00",x"28",x"55",x"55",x"04",x"24",x"55",x"55",x"00",x"00",x"00",x"00",x"00",x"04",x"28",x"28",x"00",x"00",x"00",x"00",x"2d",x"55",x"28",x"04",x"55",x"55",x"04",x"00",x"28",x"28",x"04",x"00",x"28",x"28",x"04",x"00",x"51",x"55",x"29",x"28",x"55",x"51",x"00",x"2d",x"55",x"55",x"2d",x"04",x"51",x"35",x"28",x"00",x"55",x"55",x"28",x"04",x"55",x"31",x"00",x"4d",x"55",x"04",x"28",x"55",x"55",x"04",x"24",x"55",x"55",x"28",x"00",x"51",x"55",x"04",x"28",x"55",x"28",x"00",x"51",x"51",x"00",x"2c",x"55",x"51",x"00",x"08",x"28",x"00",x"04",x"55",x"51",x"00",x"04",x"28",x"28",x"00",x"31",x"55",x"2d",x"00",x"51",x"55",x"28",x"08",x"55",x"28",x"04",x"55",x"55",x"28",x"28",x"55",x"55",x"00",x"04",x"55",x"55",x"29",x"04",x"55",x"55",x"28",x"00",x"28",x"28",x"04",x"04",x"55",x"31",x"00",x"28",x"00",x"2d",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"28",x"55",x"51",x"00",x"28",x"55",x"55",x"2d",x"00",x"31",x"35",x"31",x"00",x"28",x"55",x"35",x"2d",x"00",x"2d",x"55",x"2d",x"00",x"28",x"28",x"08",x"00",x"51",x"51",x"00",x"2d",x"2d",x"00",x"51",x"51",x"00",x"28",x"55",x"29",x"00",x"08",x"28",x"00",x"04",x"2c",x"08",x"00",x"4d",x"51",x"00",x"28",x"51",x"00",x"04",x"28",x"00",x"28",x"51",x"00",x"04",x"08",x"00",x"51",x"29",x"00",x"28",x"04",x"00",x"51",x"51",x"28",x"55",x"51",x"00",x"51",x"55",x"51",x"04",x"51",x"55",x"28",x"00",x"28",x"28",x"28",x"00",x"31",x"55",x"28",x"00",x"28",x"28",x"00",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"0c",x"04",x"55",x"51",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"55",x"35",x"2d",x"28",x"55",x"55",x"2d",x"00",x"2d",x"35",x"31",x"00",x"24",x"55",x"04",x"28",x"55",x"2d",x"00",x"51"),
(x"51",x"55",x"00",x"2c",x"35",x"31",x"04",x"31",x"35",x"2c",x"00",x"2d",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"55",x"55",x"04",x"2d",x"55",x"4d",x"00",x"4d",x"55",x"2d",x"00",x"31",x"35",x"04",x"00",x"55",x"2d",x"00",x"4d",x"55",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2d",x"04",x"51",x"55",x"28",x"00",x"31",x"35",x"2d",x"00",x"4d",x"55",x"51",x"00",x"28",x"55",x"51",x"00",x"2c",x"35",x"31",x"00",x"31",x"51",x"00",x"28",x"55",x"28",x"00",x"35",x"35",x"04",x"04",x"55",x"31",x"00",x"28",x"35",x"31",x"00",x"51",x"55",x"04",x"28",x"55",x"28",x"00",x"55",x"31",x"00",x"2c",x"35",x"04",x"04",x"55",x"28",x"00",x"31",x"2d",x"00",x"2d",x"31",x"00",x"31",x"2d",x"00",x"2d",x"31",x"00",x"51",x"2d",x"04",x"55",x"04",x"00",x"35",x"04",x"28",x"2d",x"00",x"51",x"04",x"28",x"28",x"00",x"2d",x"00",x"2d",x"2c",x"00",x"4d",x"00",x"08",x"55",x"04",x"04",x"55",x"04",x"08",x"55",x"04",x"08",x"35",x"08",x"04",x"55",x"2c",x"00",x"51",x"04",x"04",x"51",x"04",x"2c",x"35",x"04",x"04",x"55",x"28",x"04",x"55",x"04",x"04",x"51",x"00",x"2c",x"31",x"00",x"51",x"29",x"00",x"4d",x"00",x"2d",x"04",x"04",x"31",x"00",x"28",x"35",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"28",x"55",x"29",x"00",x"51",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"28",x"35",x"04",x"04",x"55",x"28",x"00",x"51",x"51",x"00",x"2c",x"31",x"00",x"2d",x"31",x"00",x"31",x"51",x"00",x"2d",x"51",x"00",x"2c",x"35",x"00",x"28",x"55",x"00",x"24",x"51",x"00",x"28",x"55",x"00",x"28",x"51",x"00",x"29",x"29",x"00",x"51",x"28",x"04",x"31",x"00",x"2d",x"04",x"04",x"51",x"00",x"31",x"08",x"04",x"51",x"00",x"29",x"2d",x"00",x"51",x"04",x"28",x"2d",x"00",x"2d",x"04",x"31",x"04",x"31",x"2c",x"00",x"51",x"28",x"00",x"55",x"04",x"28",x"35",x"04",x"08",x"35",x"08",x"00",x"51",x"2d",x"00",x"51",x"4d",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"28",x"2c",x"04",x"04",x"35",x"55",x"04",x"2c",x"35",x"31",x"00",x"28",x"55",x"31",x"00",x"4d",x"75",x"28",x"00",x"51",x"55",x"28",x"04",x"2c",x"28",x"00",x"04",x"2c",x"28",x"00",x"2d",x"35",x"2c",x"00",x"51",x"51",x"00",x"04",x"2c",x"04",x"04",x"35",x"55",x"04",x"04",x"55",x"51",x"00",x"28",x"2c",x"28",x"00",x"2d",x"55",x"51",x"00",x"28",x"2c",x"04",x"2d",x"35",x"08",x"04",x"35",x"35",x"04",x"24",x"55",x"55",x"2d",x"00",x"51",x"55",x"29",x"00",x"31",x"35",x"28",x"28",x"35",x"51",x"00",x"2c",x"35",x"35",x"2c",x"04",x"35",x"35",x"28",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"2d",x"35",x"04",x"08",x"35",x"35",x"04",x"04",x"35",x"55",x"28",x"00",x"31",x"35",x"04",x"28",x"35",x"28",x"00",x"51",x"31",x"00",x"2c",x"35",x"31",x"00",x"51",x"55",x"04",x"04",x"35",x"31",x"00",x"4d",x"55",x"4d",x"00",x"31",x"35",x"2c",x"00",x"31",x"55",x"28",x"08",x"35",x"28",x"04",x"55",x"35",x"28",x"28",x"35",x"35",x"04",x"04",x"55",x"35",x"28",x"04",x"35",x"35",x"28",x"24",x"55",x"55",x"29",x"04",x"35",x"31",x"00",x"4d",x"00",x"31",x"35",x"2c",x"00",x"28",x"2c",x"2c",x"00",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"28",x"35",x"31",x"00",x"28",x"35",x"35",x"2d",x"00",x"31",x"35",x"31",x"00",x"28",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"51",x"55",x"4d",x"00",x"31",x"51",x"00",x"2d",x"2d",x"00",x"31",x"31",x"00",x"28",x"55",x"28",x"00",x"51",x"51",x"00",x"28",x"55",x"51",x"00",x"2d",x"55",x"00",x"08",x"31",x"00",x"28",x"51",x"00",x"28",x"51",x"00",x"4d",x"4d",x"00",x"31",x"28",x"00",x"51",x"2d",x"00",x"31",x"31",x"28",x"35",x"31",x"04",x"31",x"35",x"51",x"04",x"31",x"35",x"28",x"00",x"51",x"55",x"4d",x"00",x"31",x"35",x"28",x"00",x"55",x"55",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"04",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"0c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"28",x"35",x"35",x"2d",x"00",x"2d",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"51"),
(x"55",x"35",x"04",x"2c",x"35",x"31",x"04",x"31",x"35",x"2c",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"55",x"2d",x"00",x"2d",x"55",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2d",x"00",x"2d",x"55",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"31",x"35",x"28",x"00",x"31",x"35",x"2c",x"00",x"2d",x"35",x"51",x"00",x"28",x"55",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"28",x"55",x"28",x"04",x"35",x"35",x"04",x"04",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"31",x"55",x"04",x"28",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"04",x"04",x"55",x"28",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"04",x"35",x"04",x"00",x"35",x"04",x"28",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"2d",x"00",x"2d",x"2c",x"00",x"4d",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"08",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"55",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"28",x"00",x"31",x"00",x"2d",x"08",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"28",x"55",x"28",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"28",x"35",x"04",x"04",x"35",x"28",x"00",x"51",x"31",x"00",x"2c",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"2c",x"35",x"00",x"28",x"35",x"00",x"04",x"51",x"00",x"28",x"35",x"04",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"28",x"2c",x"00",x"31",x"04",x"08",x"2d",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"28",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2d",x"00",x"51",x"2d",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2d",x"55",x"28",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"28",x"35",x"31",x"00",x"2d",x"55",x"28",x"00",x"31",x"35",x"28",x"28",x"55",x"51",x"00",x"24",x"55",x"51",x"00",x"2c",x"35",x"2c",x"00",x"31",x"51",x"00",x"28",x"55",x"28",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"51",x"55",x"4d",x"00",x"2d",x"35",x"31",x"00",x"51",x"55",x"24",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"55",x"35",x"2c",x"00",x"51",x"55",x"28",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"28",x"00",x"31",x"35",x"04",x"28",x"35",x"08",x"00",x"31",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"55",x"04",x"04",x"35",x"31",x"00",x"2c",x"55",x"2d",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"28",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"55",x"55",x"28",x"04",x"35",x"31",x"00",x"4d",x"00",x"31",x"15",x"2c",x"00",x"4d",x"55",x"55",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"28",x"35",x"35",x"2d",x"00",x"31",x"35",x"35",x"00",x"28",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"08",x"35",x"2c",x"00",x"31",x"51",x"00",x"28",x"55",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"28",x"51",x"00",x"08",x"31",x"00",x"2d",x"31",x"00",x"31",x"28",x"00",x"51",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"31",x"04",x"31",x"35",x"28",x"00",x"51",x"35",x"2d",x"00",x"31",x"35",x"08",x"00",x"55",x"55",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"04",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"0c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"2d",x"00",x"2d",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"04",x"31",x"35",x"2d",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2d",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2d",x"35",x"04",x"2c",x"15",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"28",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"28",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"28",x"04",x"35",x"35",x"04",x"04",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"28",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"04",x"04",x"35",x"28",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"04",x"31",x"00",x"2d",x"2c",x"00",x"2d",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"08",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"31",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"35",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"28",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2d",x"35",x"00",x"2c",x"35",x"00",x"28",x"35",x"00",x"04",x"31",x"00",x"2c",x"35",x"04",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"28",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"31",x"00",x"2d",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"28",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"28",x"08",x"35",x"31",x"00",x"24",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"31",x"00",x"08",x"35",x"28",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"00",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"28",x"00",x"31",x"35",x"04",x"28",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"2d",x"00",x"31",x"35",x"2c",x"00",x"2d",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"28",x"35",x"35",x"2d",x"00",x"31",x"35",x"35",x"00",x"28",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"28",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"28",x"35",x"00",x"08",x"31",x"00",x"2c",x"31",x"00",x"31",x"28",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"28",x"00",x"31",x"35",x"2d",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"04",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"0c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"15",x"2d",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2d",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"30",x"00",x"2c",x"35",x"04",x"2c",x"15",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"31",x"2c",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"31",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"35",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"30",x"31",x"00",x"31",x"31",x"00",x"2d",x"35",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"04",x"31",x"00",x"0c",x"35",x"04",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"2d",x"00",x"30",x"31",x"00",x"31",x"31",x"00",x"2d",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"28",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"28",x"08",x"35",x"35",x"00",x"04",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"28",x"08",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"15",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"28",x"35",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"35",x"35",x"00",x"30",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"28",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"28",x"35",x"00",x"08",x"31",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"00",x"31",x"15",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2d",x"08",x"35",x"15",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2d",x"00",x"30",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"30",x"00",x"30",x"35",x"04",x"2c",x"15",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"15",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"31",x"2c",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"35",x"04",x"04",x"35",x"00",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"31",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"35",x"00",x"31",x"35",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2d",x"35",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"04",x"31",x"00",x"0c",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"30",x"31",x"00",x"31",x"31",x"00",x"2d",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"28",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"35",x"35",x"00",x"30",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"00",x"31",x"15",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"04",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2d",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2d",x"00",x"30",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"30",x"35",x"04",x"2c",x"15",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"31",x"2c",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"04",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"00",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"31",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"35",x"00",x"31",x"35",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2d",x"35",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"04",x"31",x"00",x"0c",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"30",x"31",x"00",x"31",x"31",x"00",x"2d",x"35",x"08",x"04",x"35",x"35",x"04",x"0c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"28",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"30",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"35",x"35",x"00",x"30",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"00",x"31",x"15",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"04",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2d",x"08",x"35",x"35",x"30",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2d",x"00",x"30",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"30",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"30",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"31",x"2c",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"04",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"31",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"35",x"00",x"31",x"35",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2d",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"0c",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"30",x"31",x"00",x"31",x"31",x"00",x"2d",x"35",x"08",x"04",x"35",x"35",x"04",x"0c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"0c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"30",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"28",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"28",x"35",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"30",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"00",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2d",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2d",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"30",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"04",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"31",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"35",x"00",x"31",x"35",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2d",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2d",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"0c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"28",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"0c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"28",x"35",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"31",x"00",x"31",x"28",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2d",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2d",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"30",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"28",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"31",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"04",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"0c",x"35",x"04",x"04",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"31",x"00",x"2c",x"08",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"35",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"28",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"28",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"28",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"0c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"28",x"35",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"31",x"00",x"31",x"28",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2d",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2d",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2d",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"30",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"31",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"04",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"31",x"00",x"2c",x"08",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"35",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"28",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"08",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"28",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"28",x"35",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"31",x"00",x"31",x"28",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"0c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"04",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"31",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"28",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"28",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"31",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"31",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"31",x"00",x"31",x"28",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"31",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"31",x"00",x"31",x"28",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"31",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"31",x"00",x"31",x"28",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"31",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"31",x"00",x"31",x"28",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"31",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"2d",x"00",x"51",x"28",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"31",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2d",x"4d",x"00",x"28",x"04",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"31",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2d",x"4d",x"00",x"00",x"00",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"2d",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"31",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"4d",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"51",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"08",x"35",x"00",x"28",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"35",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"2d",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"04",x"2d",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"28",x"35",x"00",x"04",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"55",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"04",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"00",x"04",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"31",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"28",x"35",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"31",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"2c",x"55",x"04",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"00",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"0c",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"51",x"2c",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"28",x"55",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"24",x"2d",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"00",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"2c",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"28",x"24",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"00",x"04",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"04",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"00",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"2c",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"00",x"31",x"00",x"2d",x"04",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"00",x"00",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"28",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"31",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"08",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"2c",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"00",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2c",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"0c",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"00",x"00",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"28",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"31",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"00",x"28",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"2d",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"00",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"0c",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"00",x"00",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"51",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"55",x"00",x"24",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"04",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"51",x"51",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"00",x"00",x"2c",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"08",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"2d",x"04",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"00",x"00",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"51",x"51",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"31",x"00",x"2d",x"51",x"00",x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"4d",x"51",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"30",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"31",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"00",x"00",x"2d",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2d",x"51",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"28",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"04",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"00",x"00",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"04",x"04",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"28",x"35",x"31",x"00",x"29",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"04",x"04",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"30",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"51",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"00",x"00",x"2d",x"24",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"2d",x"2d",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"28",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"00",x"00",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"28",x"35",x"31",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"30",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"04",x"51",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"00",x"00",x"2d",x"24",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"04",x"04",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"28",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"00",x"00",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"28",x"35",x"08",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"28",x"55",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"30",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"2d",x"00",x"2c",x"31",x"00",x"31",x"0c",x"00",x"00",x"00",x"28",x"04",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"28",x"35",x"00",x"08",x"31",x"00",x"2c",x"2c",x"00",x"31",x"08",x"04",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"31",x"04",x"00",x"00",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"28",x"55",x"28",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"24",x"31",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"04",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"2c",x"35",x"00",x"08",x"31",x"00",x"28",x"28",x"00",x"31",x"08",x"04",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"04",x"51",x"00",x"00",x"00",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"28",x"55",x"28",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"31",x"2c",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"00",x"04",x"31",x"00",x"0c",x"35",x"00",x"08",x"31",x"00",x"29",x"29",x"00",x"31",x"08",x"04",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"00",x"51",x"00",x"00",x"00",x"00",x"35",x"08",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"04",x"2d",x"04",x"00",x"00",x"00",x"00",x"2d",x"55",x"51",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"31",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"51",x"29",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"04",x"51",x"00",x"0c",x"35",x"00",x"08",x"31",x"00",x"04",x"04",x"00",x"31",x"08",x"00",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"00",x"28",x"00",x"00",x"00",x"00",x"51",x"28",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"04",x"2c",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"2d",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"24",x"51",x"00",x"0c",x"35",x"00",x"08",x"31",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"28",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"31",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"51",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"2d",x"31",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"08",x"00",x"2c",x"35",x"00",x"08",x"31",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"51",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"2d",x"2d",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"31",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"2c",x"35",x"00",x"08",x"31",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"4d",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"04",x"04",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"04",x"08",x"28",x"00",x"2d",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"0c",x"35",x"00",x"08",x"31",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"55",x"51",x"00",x"2c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"2d",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"35",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"0c",x"35",x"00",x"08",x"31",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"31",x"31",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"51",x"2d",x"00",x"2c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"2d",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"55",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2d",x"31",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"0c",x"35",x"00",x"08",x"31",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"31",x"2c",x"00",x"51",x"51",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"35"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"08",x"00",x"04",x"00",x"00",x"2c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"4d",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"08",x"35",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"51",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"2d",x"51",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"0c",x"35",x"00",x"08",x"31",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"30",x"35",x"04",x"08",x"35",x"35",x"04",x"08",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"2d",x"2d",x"00",x"28",x"2d",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"51"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"28",x"00",x"00",x"00",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"28",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"08",x"55",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"04",x"51",x"04",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"28",x"2c",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"0c",x"35",x"00",x"08",x"31",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"30",x"35",x"04",x"08",x"35",x"35",x"04",x"04",x"35",x"35",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"55",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"35",x"35",x"00",x"2d",x"2d",x"00",x"00",x"00",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"51"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"28",x"00",x"00",x"00",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"00",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"04",x"28",x"55",x"04",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"2d",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"0c",x"35",x"00",x"28",x"31",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"30",x"35",x"04",x"08",x"35",x"35",x"04",x"24",x"55",x"55",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"55",x"04",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"35",x"35",x"00",x"2d",x"2d",x"00",x"00",x"00",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"2c"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2d",x"35",x"31",x"00",x"00",x"00",x"00",x"28",x"55",x"28",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"08",x"35",x"28",x"00",x"00",x"00",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"00",x"00",x"2c",x"2c",x"00",x"31",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"04",x"28",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"51",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"0c",x"35",x"00",x"28",x"51",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"28",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"31",x"31",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"30",x"35",x"04",x"08",x"35",x"35",x"04",x"24",x"55",x"55",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"28",x"00",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"4d",x"2d",x"00",x"00",x"00",x"00",x"28",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2d",x"55",x"51",x"00",x"00",x"00",x"00",x"28",x"55",x"28",x"00",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"28",x"35",x"28",x"00",x"00",x"00",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"00",x"00",x"2c",x"2c",x"00",x"2d",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"51",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"0c",x"35",x"00",x"28",x"51",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"28",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"2d",x"51",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"30",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"28",x"28",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"28",x"55",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"04",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"08",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"28",x"35",x"28",x"00",x"00",x"00",x"00",x"0c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"00",x"00",x"2c",x"2c",x"00",x"51",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"0c",x"35",x"04",x"00",x"04",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"28",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"4d",x"51",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"24",x"55",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"75",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"39",x"2c",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"08",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"28",x"55",x"28",x"00",x"00",x"00",x"00",x"2c",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"2d",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"08",x"28",x"00",x"00",x"00",x"2c",x"2c",x"00",x"4d",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"04",x"04",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2d",x"55",x"28",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"24",x"51",x"51",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"51",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"08",x"35",x"2c",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"35",x"35",x"28",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"28",x"55",x"28",x"00",x"00",x"00",x"00",x"2c",x"35",x"04",x"04",x"35",x"08",x"00",x"31",x"2d",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"28",x"28",x"00",x"00",x"00",x"2c",x"2c",x"00",x"04",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"2d",x"51",x"24",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"31",x"35",x"04",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"51",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"28",x"35",x"2c",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"31",x"35",x"28",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"04",x"04",x"35",x"08",x"00",x"51",x"2d",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"28",x"28",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"08",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"04",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"2d",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"04",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"28",x"55",x"2d",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"04",x"55",x"55",x"28",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"55",x"04",x"04",x"35",x"08",x"00",x"4d",x"29",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"28",x"28",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"55",x"28",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"55",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"4d",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"24",x"51",x"28",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"51",x"55",x"28",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"55",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"28",x"28",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"55",x"28",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"04",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"31",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"2c",x"4d",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"2d",x"2d",x"24",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"2d",x"00",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"04",x"24",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"2d",x"04",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0c",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"00",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"2d",x"55",x"2d",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"55",x"31",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"55",x"51",x"00",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"28",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0c",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"51",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"28",x"2c",x"28",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"51",x"51",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"51",x"55",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"2c",x"28",x"00",x"31",x"15",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"24",x"55",x"04",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"28",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"28",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"51",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"31",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"28",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"28",x"28",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"24",x"55",x"04",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"28",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4d",x"51",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"28",x"35",x"04",x"00",x"00",x"00",x"28",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"51",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"51",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"0c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"55",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"35",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"00",x"28",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"28",x"35",x"04",x"00",x"00",x"00",x"28",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"4d",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"4d",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"0c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"04",x"51",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"31",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"28",x"35",x"04",x"00",x"00",x"00",x"28",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"0c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"15",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"55",x"08",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"51",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"28",x"35",x"04",x"00",x"00",x"00",x"28",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"31",x"04",x"08",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"51",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"51",x"28",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"51",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"2d",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"28",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"31",x"04",x"28",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"35",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"15",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2d",x"2d",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"51",x"28",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"2d",x"04",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"51",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"0c",x"35",x"04",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"31",x"04",x"28",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"04",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"00",x"35",x"35",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"51",x"24",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"31",x"04",x"28",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"2d",x"55",x"04",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"00",x"55",x"35",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"55",x"2d",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"35",x"04",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"51",x"51",x"04",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"28",x"04",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"28",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"31",x"04",x"04",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"4d",x"51",x"24",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"00",x"51",x"55",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"55",x"4d",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"55",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"28",x"55",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"28",x"00",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"28",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"28",x"28",x"04",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"00",x"28",x"28",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"2c",x"28",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"51",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"51",x"51",x"04",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"28",x"51",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"55",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"28",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2d",x"55",x"2d",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4d",x"51",x"51",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"04",x"08",x"00",x"00",x"35",x"2c",x"00",x"2c",x"35",x"04",x"2d",x"55",x"51",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"00",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"51",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"2c",x"51",x"28",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"08",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"28",x"31",x"2d",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2c",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"35",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"2c",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"55",x"04",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"04",x"04",x"04",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"55",x"35",x"04",x"04",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"04",x"31",x"35",x"2d",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"04",x"04",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"04",x"55",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"2d",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"51",x"00",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"31",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"08",x"04",x"31",x"2d",x"00",x"04",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"30",x"00",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"04",x"31",x"35",x"2d",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"31",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"00",x"4d",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"28",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"51",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"04",x"04",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"30",x"00",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"04",x"31",x"35",x"2d",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"2d",x"51",x"00",x"2c",x"35",x"00",x"08",x"35",x"04",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"35",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"51",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"31",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2d",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"51",x"55",x"4d",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"2c",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"08",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"28",x"28",x"00",x"2c",x"35",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"31",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"28",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"2c",x"35",x"51",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"4d",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2d",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"28",x"2c",x"24",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"08",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"2d",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"04",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"51",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"51",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"28",x"55",x"51",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"28",x"2c",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2d",x"55",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"28",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"55",x"04",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"51",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"51",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"04",x"28",x"28",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"55",x"2d",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"08",x"35",x"35",x"31",x"00",x"2d",x"51",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"28",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"51",x"04",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"28",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"28",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"51",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"28",x"35",x"35",x"2d",x"00",x"04",x"28",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"08",x"00",x"35",x"04",x"28",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"28",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"28",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"04",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"28",x"35",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"55",x"51",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"08",x"00",x"35",x"04",x"28",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"55",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"28",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"28",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"28",x"55",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"51",x"2d",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"24",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"55",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"28",x"55",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"28",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"04",x"35",x"35",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2c",x"24",x"31",x"31",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"35",x"04",x"00",x"35",x"04",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"2d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"24",x"2d",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"00",x"35",x"35",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"2d",x"00",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"55",x"04",x"00",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"00",x"51",x"55",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"28",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"04",x"55",x"24",x"00",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"0c",x"00",x"2c",x"2c",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"28",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"2d",x"00",x"31",x"31",x"00",x"35",x"2c",x"00",x"28",x"00",x"00",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"28",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"08",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"2d",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"04",x"00",x"31",x"31",x"00",x"35",x"30",x"00",x"00",x"00",x"04",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"08",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4d",x"55",x"28",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"28",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"4d",x"51",x"51",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"35",x"31",x"00",x"00",x"00",x"04",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"55",x"28",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"00",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"28",x"55",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"55",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"04",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"55",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"35",x"31",x"00",x"00",x"00",x"04",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"51",x"24",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"28",x"51",x"51",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"04",x"51",x"51",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"51",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"35",x"31",x"00",x"00",x"00",x"04",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"00",x"04",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"00",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"35",x"31",x"00",x"00",x"00",x"04",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"15",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"35",x"31",x"00",x"00",x"00",x"04",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"55",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"35",x"31",x"00",x"00",x"00",x"04",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"2d",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"0c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"35",x"31",x"00",x"00",x"00",x"04",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"51",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"2c",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"35",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"35",x"31",x"00",x"00",x"00",x"04",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"51",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2c",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"28",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"31",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"51",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"51",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"35",x"31",x"00",x"00",x"00",x"04",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"28",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2d",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2d",x"55",x"55",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"55",x"28",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"51",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"04",x"51",x"55",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"51",x"55",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"35",x"31",x"00",x"00",x"00",x"04",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2d",x"55",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"2d",x"55",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"04",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"51",x"55",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"15",x"31",x"00",x"08",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"31",x"00",x"35",x"31",x"00",x"00",x"00",x"04",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"2d",x"55",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"04",x"08",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"04",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"31",x"00",x"35",x"31",x"00",x"00",x"00",x"00",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"51",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"55",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4d",x"4d",x"00",x"35",x"31",x"00",x"00",x"00",x"00",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"55",x"55",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"2c",x"55",x"51",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2c",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"4d",x"00",x"35",x"31",x"00",x"00",x"00",x"00",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"51",x"04",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"2d",x"55",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"28",x"51",x"2d",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2d",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"31",x"00",x"00",x"00",x"00",x"4d",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2c",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"55",x"55",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"28",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"28",x"51",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"2d",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"0c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2d",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"04",x"4d",x"4d",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"28",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2d",x"00",x"2d",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"2c",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"2d",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"04",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"08",x"35",x"28",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"28",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"35",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"4d",x"55",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"28",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"04",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"28",x"55",x"28",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"28",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"55",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"04",x"28",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"55",x"28",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"28",x"55",x"28",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"08",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"08",x"35",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4d",x"55",x"28",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2c",x"35",x"31",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"55",x"28",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"55",x"31",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"08",x"35",x"35",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"08",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"51",x"55",x"28",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"28",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"2d",x"55",x"2d",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"51",x"4d",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"04",x"35",x"31",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"51",x"51",x"24",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"28",x"55",x"55",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"29",x"51",x"2d",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"24",x"55",x"51",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"08",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"28",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"28",x"51",x"51",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"04",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"24",x"51",x"51",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"28",x"35",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"55",x"28",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4d",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"28",x"00",x"04",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"28",x"35",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"31",x"24",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"35",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"28",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"28",x"55",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"08",x"35",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"35",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"28",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"24",x"2d",x"2d",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"04",x"51",x"55",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"55",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"04",x"2c",x"2c",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"28",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"08",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"28",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"08",x"00",x"31",x"35",x"0c",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"0c",x"28",x"55",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"55",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"28",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"24",x"51",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"51",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"28",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"55",x"51",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"28",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"51",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"0c",x"04",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"15",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"35",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"0c",x"04",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"08",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"0c",x"04",x"55",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"0c",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"35",x"35",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"0c",x"24",x"55",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"55",x"51",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"0c",x"00",x"2c",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"0c",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"2c",x"28",x"00",x"04",x"35",x"35",x"0c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"28",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"08",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"28",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"28",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"28",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"28",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"28",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"51",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"28",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"35",x"55",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"28",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"28",x"2d",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"28",x"35",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"04",x"04",x"55",x"55",x"04",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"31",x"35",x"28",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"28",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"28",x"55",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"55",x"04",x"00",x"28",x"28",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"28",x"00",x"51",x"55",x"28",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"55",x"35",x"2c",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"55",x"55",x"28",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"04",x"28",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"51",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"55",x"28",x"00",x"08",x"08",x"04",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"51",x"51",x"29",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"51",x"55",x"28",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"51",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"04",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"04",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"0c",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"15",x"0c",x"04",x"55",x"55",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"2c",x"00",x"51",x"51",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"08",x"35",x"35",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2c",x"00",x"31",x"35",x"2c",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"35",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"28",x"55",x"35",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2d",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"55",x"31",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"28",x"55",x"55",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2d",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"04",x"55",x"51",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"04",x"2c",x"28",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2d",x"00",x"51",x"55",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2c",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"00",x"08",x"04",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"35",x"35",x"04",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2d",x"00",x"08",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"31",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"08",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"55",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"51",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"51",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"28",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"04",x"51",x"51",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"2d",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"55",x"55",x"28",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"30",x"35",x"35",x"04",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"0c",x"00",x"35",x"35",x"04",x"08",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"31",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"51",x"51",x"24",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"28",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"51",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"55",x"51",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"15",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"24",x"51",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"2d",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"31",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"31",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2d",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"4d",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"55",x"2d",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"28",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"4d",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"55",x"4d",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"04",x"00",x"31",x"35",x"2c",x"00",x"31",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08",x"04",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"2d",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"2d",x"55",x"55",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"4d",x"51",x"51",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"51",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"55",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"4d",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"2d",x"2d",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"08",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"28",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"28",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"28",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"28",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"08",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"28",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"35",x"28",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"28",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2d",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"55",x"28",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"04",x"2d",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4d",x"55",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4d",x"55",x"28",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"2c",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"2c",x"04",x"00",x"35",x"35",x"04",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"31",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"51",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"28",x"2d",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"55",x"55",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"51",x"51",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"2c",x"2c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"35",x"35",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"51",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")


);
	



-- one bit mask  0 - off 1 dispaly 
type object_form is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object : object_form := (

("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111")
);





signal bCoord_X : integer := 0;-- offset from start position 
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';

--		
signal objectEndX : integer;
signal objectEndY : integer;

begin

-- Calculate object end boundaries
objectEndX	<= object_X_size+ObjectStartX;
objectEndY	<= object_Y_size+ObjectStartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

-- test if ooCoord is in the rectangle defined by Start and End 
	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectEndX) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectEndY) else '0';

-- calculate offset from start corner 
	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 


process ( RESETn, CLK)

  		
   begin
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;

		elsif rising_edge(CLK) then
		
			mVGA_RGB	<=  object_colors(bCoord_Y , bCoord_X);	--get from colors table 
			drawing_request	<= object(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table if inside rectangle  
	end if;

  end process;

		
end behav;		