--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity Coin_Sound is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ENA                   : in std_logic;
  ADDR    					: in std_logic_vector(14 downto 0);
  Q       					: out std_logic_vector(15 downto 0);
  Done                  : out std_logic

  
);
end Coin_Sound;

architecture arch of Coin_Sound is
constant array_size 			: integer := 6294 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal sin_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
  sintable_proc: process(resetN, CLK)
    constant sin_table : table_type := (
---start 0 v


X"0000",
X"0000",
X"007D",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"FE89",
X"FE89",
X"0659",
X"04E2",
X"0659",
X"0177",
X"F92A",
X"FB9B",
X"FA24",
X"FF06",
X"06D6",
X"03E8",
X"05DC",
X"01F4",
X"FA24",
X"FB1E",
X"F9A7",
X"FB1E",
X"0465",
X"05DC",
X"05DC",
X"04E2",
X"FB1E",
X"FAA1",
X"FA24",
X"FB1E",
X"04E2",
X"055F",
X"05DC",
X"04E2",
X"FB1E",
X"FA24",
X"FAA1",
X"FC18",
X"055F",
X"055F",
X"04E2",
X"03E8",
X"FAA1",
X"FB1E",
X"FA24",
X"FC18",
X"055F",
X"055F",
X"055F",
X"0465",
X"FB1E",
X"F9A7",
X"FAA1",
X"FA24",
X"0271",
X"06D6",
X"04E2",
X"05DC",
X"FE0C",
X"F92A",
X"FB1E",
X"F9A7",
X"0271",
X"0659",
X"04E2",
X"05DC",
X"FD12",
X"F9A7",
X"FB1E",
X"F9A7",
X"0271",
X"0659",
X"04E2",
X"05DC",
X"FD12",
X"F92A",
X"FB1E",
X"FA24",
X"02EE",
X"06D6",
X"04E2",
X"0659",
X"00FA",
X"F92A",
X"FB9B",
X"FA24",
X"FF06",
X"06D6",
X"0465",
X"0659",
X"00FA",
X"F9A7",
X"FB1E",
X"F9A7",
X"FF06",
X"0659",
X"04E2",
X"06D6",
X"007D",
X"F92A",
X"FB9B",
X"F9A7",
X"FF83",
X"0659",
X"0465",
X"0659",
X"0000",
X"F9A7",
X"FB9B",
X"FAA1",
X"FC18",
X"04E2",
X"04E2",
X"055F",
X"03E8",
X"FAA1",
X"FB1E",
X"FA24",
X"FC18",
X"055F",
X"055F",
X"05DC",
X"036B",
X"FAA1",
X"FAA1",
X"F9A7",
X"FC95",
X"05DC",
X"055F",
X"0659",
X"036B",
X"FA24",
X"FAA1",
X"F9A7",
X"FC95",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"FC95",
X"F9A7",
X"FAA1",
X"FA24",
X"036B",
X"05DC",
X"04E2",
X"055F",
X"FC18",
X"FAA1",
X"FB1E",
X"FAA1",
X"036B",
X"055F",
X"04E2",
X"05DC",
X"FC95",
X"FA24",
X"FB1E",
X"FA24",
X"036B",
X"05DC",
X"0465",
X"05DC",
X"FC95",
X"FAA1",
X"FB1E",
X"FA24",
X"02EE",
X"05DC",
X"04E2",
X"06D6",
X"0000",
X"F9A7",
X"FB9B",
X"F9A7",
X"007D",
X"0659",
X"0465",
X"0659",
X"FF83",
X"F9A7",
X"FB1E",
X"F92A",
X"007D",
X"06D6",
X"0465",
X"0659",
X"FF06",
X"F92A",
X"FC18",
X"F9A7",
X"00FA",
X"05DC",
X"0465",
X"0659",
X"FF06",
X"F9A7",
X"FB1E",
X"FA24",
X"FD8F",
X"055F",
X"04E2",
X"05DC",
X"0271",
X"FA24",
X"FB1E",
X"FA24",
X"FD8F",
X"0659",
X"04E2",
X"05DC",
X"0271",
X"FA24",
X"FB9B",
X"FA24",
X"FD8F",
X"0659",
X"04E2",
X"05DC",
X"0271",
X"FAA1",
X"FB9B",
X"FA24",
X"FE0C",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"FC18",
X"FAA1",
X"FB1E",
X"FAA1",
X"03E8",
X"05DC",
X"04E2",
X"04E2",
X"FC18",
X"FAA1",
X"FB1E",
X"FB1E",
X"036B",
X"05DC",
X"04E2",
X"04E2",
X"FC18",
X"FA24",
X"FB1E",
X"FB1E",
X"0465",
X"05DC",
X"04E2",
X"04E2",
X"FB9B",
X"FA24",
X"FB1E",
X"FA24",
X"00FA",
X"05DC",
X"0465",
X"0659",
X"FF06",
X"F9A7",
X"FB9B",
X"F9A7",
X"0177",
X"05DC",
X"0465",
X"0659",
X"FF06",
X"FA24",
X"FB9B",
X"F9A7",
X"0177",
X"0659",
X"0465",
X"0659",
X"FE89",
X"F9A7",
X"FC18",
X"F9A7",
X"0177",
X"0659",
X"0465",
X"0659",
X"FE89",
X"F9A7",
X"FB1E",
X"F9A7",
X"FD8F",
X"0659",
X"0465",
X"0659",
X"01F4",
X"F9A7",
X"FB9B",
X"F9A7",
X"FE0C",
X"0659",
X"0465",
X"06D6",
X"01F4",
X"F9A7",
X"FB1E",
X"F9A7",
X"FE89",
X"0659",
X"0465",
X"06D6",
X"0177",
X"F92A",
X"FB9B",
X"F92A",
X"FF06",
X"0659",
X"04E2",
X"05DC",
X"0465",
X"FB1E",
X"FAA1",
X"FA24",
X"FB1E",
X"055F",
X"055F",
X"05DC",
X"0465",
X"FAA1",
X"FAA1",
X"FAA1",
X"FB9B",
X"04E2",
X"04E2",
X"05DC",
X"0465",
X"FAA1",
X"FAA1",
X"FA24",
X"FC18",
X"055F",
X"04E2",
X"0659",
X"03E8",
X"FAA1",
X"FAA1",
X"FB1E",
X"F9A7",
X"0271",
X"0659",
X"0465",
X"06D6",
X"FD8F",
X"F9A7",
X"FB1E",
X"F9A7",
X"0271",
X"0659",
X"04E2",
X"0659",
X"FD8F",
X"F9A7",
X"FAA1",
X"F9A7",
X"0271",
X"0659",
X"055F",
X"0659",
X"FD12",
X"F9A7",
X"FAA1",
X"F9A7",
X"02EE",
X"06D6",
X"04E2",
X"06D6",
X"007D",
X"F9A7",
X"FB1E",
X"F92A",
X"FF83",
X"06D6",
X"04E2",
X"06D6",
X"007D",
X"F9A7",
X"FB1E",
X"F8AD",
X"FF83",
X"06D6",
X"055F",
X"06D6",
X"007D",
X"F8AD",
X"FAA1",
X"F9A7",
X"0000",
X"0753",
X"055F",
X"0659",
X"0000",
X"F8AD",
X"FB1E",
X"F92A",
X"0000",
X"06D6",
X"055F",
X"0659",
X"036B",
X"F9A7",
X"FA24",
X"FA24",
X"FC95",
X"0659",
X"055F",
X"05DC",
X"036B",
X"F9A7",
X"FAA1",
X"F9A7",
X"FD12",
X"05DC",
X"055F",
X"05DC",
X"02EE",
X"FA24",
X"FAA1",
X"FA24",
X"FC95",
X"05DC",
X"055F",
X"0659",
X"02EE",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"036B",
X"06D6",
X"04E2",
X"05DC",
X"FC18",
X"F9A7",
X"FB1E",
X"FA24",
X"03E8",
X"05DC",
X"04E2",
X"055F",
X"FC95",
X"FA24",
X"FAA1",
X"FA24",
X"036B",
X"05DC",
X"055F",
X"055F",
X"FC18",
X"FA24",
X"FAA1",
X"FB1E",
X"036B",
X"05DC",
X"0465",
X"0659",
X"0000",
X"F9A7",
X"FB9B",
X"F92A",
X"0000",
X"0659",
X"04E2",
X"06D6",
X"0000",
X"F9A7",
X"FB1E",
X"F92A",
X"007D",
X"06D6",
X"04E2",
X"06D6",
X"0000",
X"F92A",
X"FAA1",
X"F92A",
X"007D",
X"0659",
X"04E2",
X"0753",
X"FF83",
X"F92A",
X"FAA1",
X"F92A",
X"FD12",
X"05DC",
X"055F",
X"0659",
X"02EE",
X"F9A7",
X"FAA1",
X"F9A7",
X"FD8F",
X"05DC",
X"04E2",
X"0659",
X"02EE",
X"FA24",
X"FB1E",
X"FA24",
X"FD8F",
X"05DC",
X"04E2",
X"05DC",
X"0271",
X"F9A7",
X"FB1E",
X"FA24",
X"FE0C",
X"05DC",
X"04E2",
X"05DC",
X"01F4",
X"FA24",
X"FB1E",
X"FAA1",
X"FB1E",
X"03E8",
X"055F",
X"04E2",
X"055F",
X"FC18",
X"FAA1",
X"FAA1",
X"FB1E",
X"03E8",
X"055F",
X"055F",
X"04E2",
X"FB9B",
X"FAA1",
X"FB1E",
X"FB9B",
X"03E8",
X"055F",
X"04E2",
X"04E2",
X"FB9B",
X"FAA1",
X"FAA1",
X"FB9B",
X"0465",
X"055F",
X"04E2",
X"05DC",
X"FE89",
X"F9A7",
X"FB9B",
X"F9A7",
X"0177",
X"0659",
X"0465",
X"055F",
X"FE0C",
X"FA24",
X"FB9B",
X"FA24",
X"01F4",
X"05DC",
X"0465",
X"05DC",
X"FE89",
X"FA24",
X"FB9B",
X"F9A7",
X"0177",
X"0659",
X"04E2",
X"05DC",
X"FE0C",
X"F9A7",
X"FB9B",
X"FA24",
X"FE89",
X"0659",
X"0465",
X"05DC",
X"0177",
X"F9A7",
X"FB9B",
X"FA24",
X"FE89",
X"06D6",
X"0465",
X"05DC",
X"00FA",
X"F9A7",
X"FB9B",
X"FA24",
X"FF06",
X"0659",
X"0465",
X"05DC",
X"0177",
X"FA24",
X"FB9B",
X"F9A7",
X"FF06",
X"05DC",
X"04E2",
X"05DC",
X"03E8",
X"FB9B",
X"FAA1",
X"FAA1",
X"FB9B",
X"04E2",
X"055F",
X"055F",
X"0465",
X"FAA1",
X"FB1E",
X"FAA1",
X"FB9B",
X"055F",
X"055F",
X"055F",
X"03E8",
X"FAA1",
X"FB1E",
X"FAA1",
X"FB9B",
X"055F",
X"04E2",
X"055F",
X"03E8",
X"FB1E",
X"FAA1",
X"FA24",
X"FC18",
X"0465",
X"05DC",
X"04E2",
X"05DC",
X"FD8F",
X"F9A7",
X"FB1E",
X"FA24",
X"02EE",
X"0659",
X"04E2",
X"05DC",
X"FD12",
X"FA24",
X"FB9B",
X"FA24",
X"02EE",
X"05DC",
X"04E2",
X"05DC",
X"FD8F",
X"F9A7",
X"FB1E",
X"FA24",
X"02EE",
X"05DC",
X"05DC",
X"055F",
X"FD12",
X"FA24",
X"FB9B",
X"FA24",
X"FF83",
X"06D6",
X"0465",
X"0659",
X"007D",
X"F9A7",
X"FB9B",
X"FA24",
X"0000",
X"05DC",
X"0465",
X"05DC",
X"0000",
X"FA24",
X"FB9B",
X"F9A7",
X"0000",
X"05DC",
X"0465",
X"0659",
X"007D",
X"F9A7",
X"FB1E",
X"F9A7",
X"007D",
X"0659",
X"04E2",
X"055F",
X"02EE",
X"FAA1",
X"FB1E",
X"FB1E",
X"FD12",
X"05DC",
X"0465",
X"055F",
X"036B",
X"FA24",
X"FB9B",
X"FAA1",
X"FC95",
X"055F",
X"0465",
X"05DC",
X"02EE",
X"FAA1",
X"FB1E",
X"FA24",
X"FD12",
X"055F",
X"04E2",
X"05DC",
X"0271",
X"FAA1",
X"FB1E",
X"FAA1",
X"FB1E",
X"036B",
X"05DC",
X"0465",
X"04E2",
X"FC95",
X"FA24",
X"FB9B",
X"FAA1",
X"03E8",
X"055F",
X"04E2",
X"04E2",
X"FC18",
X"FAA1",
X"FB9B",
X"FB1E",
X"036B",
X"055F",
X"0465",
X"04E2",
X"FC95",
X"FB1E",
X"FB1E",
X"FB1E",
X"036B",
X"055F",
X"055F",
X"04E2",
X"FC95",
X"F9A7",
X"FB9B",
X"FAA1",
X"00FA",
X"0659",
X"03E8",
X"05DC",
X"FF06",
X"FA24",
X"FB9B",
X"FA24",
X"00FA",
X"055F",
X"03E8",
X"0659",
X"FF06",
X"FAA1",
X"FC18",
X"F9A7",
X"00FA",
X"05DC",
X"0465",
X"0659",
X"FF06",
X"FA24",
X"FB9B",
X"F9A7",
X"01F4",
X"055F",
X"03E8",
X"0659",
X"01F4",
X"FAA1",
X"FC18",
X"F9A7",
X"FD8F",
X"05DC",
X"03E8",
X"05DC",
X"01F4",
X"FA24",
X"FC18",
X"F92A",
X"FE0C",
X"05DC",
X"0465",
X"0659",
X"0177",
X"F9A7",
X"FC18",
X"FA24",
X"FE89",
X"05DC",
X"036B",
X"0659",
X"0177",
X"FAA1",
X"FC18",
X"FA24",
X"FB9B",
X"03E8",
X"04E2",
X"04E2",
X"0465",
X"FB9B",
X"FB9B",
X"FAA1",
X"FB1E",
X"0465",
X"04E2",
X"05DC",
X"03E8",
X"FB9B",
X"FB1E",
X"FB1E",
X"FC18",
X"03E8",
X"0465",
X"0465",
X"04E2",
X"FC95",
X"FB1E",
X"FA24",
X"FB1E",
X"0465",
X"055F",
X"055F",
X"05DC",
X"FE0C",
X"F9A7",
X"FB9B",
X"FA24",
X"0271",
X"0659",
X"03E8",
X"055F",
X"FE0C",
X"FA24",
X"FB9B",
X"FAA1",
X"01F4",
X"055F",
X"03E8",
X"05DC",
X"FE0C",
X"F9A7",
X"FB9B",
X"FAA1",
X"0271",
X"0659",
X"0465",
X"04E2",
X"FD8F",
X"F9A7",
X"FB9B",
X"FB1E",
X"01F4",
X"05DC",
X"0465",
X"055F",
X"00FA",
X"FA24",
X"FC18",
X"FA24",
X"FE89",
X"04E2",
X"04E2",
X"06D6",
X"0177",
X"F9A7",
X"FB9B",
X"F9A7",
X"FF83",
X"0659",
X"0465",
X"055F",
X"007D",
X"FA24",
X"FC18",
X"FA24",
X"FF06",
X"05DC",
X"03E8",
X"0659",
X"007D",
X"FA24",
X"FB1E",
X"FB9B",
X"FD12",
X"04E2",
X"0465",
X"0465",
X"02EE",
X"FB1E",
X"FC18",
X"FB9B",
X"FC18",
X"0465",
X"03E8",
X"055F",
X"0465",
X"FC18",
X"FB1E",
X"F9A7",
X"FB9B",
X"0465",
X"0659",
X"05DC",
X"02EE",
X"FA24",
X"FA24",
X"FB9B",
X"FD12",
X"04E2",
X"04E2",
X"0465",
X"055F",
X"FE0C",
X"FAA1",
X"FB1E",
X"FAA1",
X"0271",
X"0659",
X"04E2",
X"04E2",
X"FC18",
X"FAA1",
X"FB1E",
X"007D",
X"05DC",
X"055F",
X"FE89",
X"FB1E",
X"FB1E",
X"0177",
X"055F",
X"055F",
X"FD12",
X"FB1E",
X"FA24",
X"0000",
X"055F",
X"055F",
X"0000",
X"FB1E",
X"FA24",
X"01F4",
X"055F",
X"05DC",
X"007D",
X"FA24",
X"FA24",
X"0000",
X"05DC",
X"05DC",
X"FF83",
X"FAA1",
X"F9A7",
X"01F4",
X"055F",
X"0659",
X"007D",
X"FA24",
X"FAA1",
X"0000",
X"05DC",
X"055F",
X"FE0C",
X"FA24",
X"FB1E",
X"0271",
X"055F",
X"05DC",
X"0000",
X"F9A7",
X"FA24",
X"01F4",
X"0659",
X"05DC",
X"FD8F",
X"F9A7",
X"FA24",
X"FF06",
X"0659",
X"05DC",
X"FF06",
X"F9A7",
X"FB1E",
X"01F4",
X"0659",
X"04E2",
X"FD12",
X"FA24",
X"FA24",
X"0000",
X"055F",
X"055F",
X"FE89",
X"FAA1",
X"FB1E",
X"01F4",
X"055F",
X"04E2",
X"007D",
X"FB1E",
X"FAA1",
X"00FA",
X"05DC",
X"04E2",
X"FE0C",
X"F92A",
X"FB1E",
X"036B",
X"05DC",
X"05DC",
X"0000",
X"FA24",
X"FAA1",
X"007D",
X"055F",
X"055F",
X"FF06",
X"FB1E",
X"FAA1",
X"FE89",
X"04E2",
X"055F",
X"007D",
X"FAA1",
X"FB1E",
X"00FA",
X"05DC",
X"055F",
X"FD8F",
X"FA24",
X"FB1E",
X"FF06",
X"05DC",
X"055F",
X"0000",
X"FAA1",
X"F9A7",
X"00FA",
X"05DC",
X"05DC",
X"0177",
X"FB1E",
X"FA24",
X"FF06",
X"055F",
X"05DC",
X"0000",
X"FAA1",
X"FAA1",
X"00FA",
X"055F",
X"055F",
X"0177",
X"FAA1",
X"FA24",
X"0000",
X"05DC",
X"05DC",
X"FF83",
X"F9A7",
X"FA24",
X"01F4",
X"055F",
X"0659",
X"0177",
X"F9A7",
X"FA24",
X"FF06",
X"05DC",
X"0659",
X"FF83",
X"FAA1",
X"FA24",
X"FD12",
X"05DC",
X"05DC",
X"00FA",
X"FAA1",
X"FA24",
X"007D",
X"0659",
X"055F",
X"FE89",
X"FA24",
X"FA24",
X"FF06",
X"05DC",
X"05DC",
X"007D",
X"F9A7",
X"F9A7",
X"007D",
X"055F",
X"05DC",
X"02EE",
X"FAA1",
X"FA24",
X"FE89",
X"055F",
X"05DC",
X"007D",
X"FA24",
X"FA24",
X"007D",
X"055F",
X"05DC",
X"01F4",
X"FAA1",
X"FA24",
X"FF06",
X"055F",
X"055F",
X"0000",
X"FAA1",
X"FAA1",
X"FC95",
X"04E2",
X"05DC",
X"01F4",
X"FB1E",
X"F9A7",
X"FF83",
X"0465",
X"05DC",
X"0000",
X"FAA1",
X"FAA1",
X"FD8F",
X"0465",
X"05DC",
X"0177",
X"FB1E",
X"FA24",
X"FF06",
X"055F",
X"055F",
X"02EE",
X"FB1E",
X"FA24",
X"FE0C",
X"04E2",
X"05DC",
X"00FA",
X"FB1E",
X"FB1E",
X"FF06",
X"055F",
X"055F",
X"036B",
X"FB1E",
X"F9A7",
X"FE0C",
X"04E2",
X"0659",
X"0177",
X"FAA1",
X"FA24",
X"FF06",
X"04E2",
X"0659",
X"0271",
X"FB1E",
X"FA24",
X"FE89",
X"04E2",
X"055F",
X"00FA",
X"FAA1",
X"FA24",
X"FC18",
X"055F",
X"0659",
X"01F4",
X"FAA1",
X"F9A7",
X"FF06",
X"055F",
X"0659",
X"007D",
X"F9A7",
X"FA24",
X"FD12",
X"055F",
X"05DC",
X"01F4",
X"FA24",
X"FA24",
X"FF06",
X"05DC",
X"0659",
X"036B",
X"FAA1",
X"FA24",
X"FE0C",
X"055F",
X"0659",
X"00FA",
X"FA24",
X"F92A",
X"FF06",
X"05DC",
X"05DC",
X"02EE",
X"FB1E",
X"FA24",
X"FE0C",
X"055F",
X"055F",
X"00FA",
X"FA24",
X"FAA1",
X"FD8F",
X"04E2",
X"055F",
X"01F4",
X"FAA1",
X"FA24",
X"FF06",
X"055F",
X"06D6",
X"007D",
X"FA24",
X"FAA1",
X"FD12",
X"04E2",
X"0659",
X"0271",
X"FB1E",
X"FA24",
X"FE89",
X"05DC",
X"055F",
X"0177",
X"FAA1",
X"FA24",
X"FD12",
X"055F",
X"05DC",
X"0177",
X"FB1E",
X"FA24",
X"FF06",
X"05DC",
X"055F",
X"036B",
X"FB9B",
X"FA24",
X"FD8F",
X"055F",
X"05DC",
X"01F4",
X"FAA1",
X"F9A7",
X"FF06",
X"055F",
X"05DC",
X"03E8",
X"FB1E",
X"FA24",
X"FD8F",
X"04E2",
X"05DC",
X"0177",
X"FAA1",
X"FAA1",
X"FC18",
X"03E8",
X"05DC",
X"02EE",
X"FB9B",
X"FA24",
X"FE0C",
X"04E2",
X"05DC",
X"00FA",
X"FAA1",
X"FAA1",
X"FC95",
X"0465",
X"05DC",
X"02EE",
X"FB9B",
X"FAA1",
X"FE0C",
X"055F",
X"04E2",
X"03E8",
X"FC95",
X"FAA1",
X"FD12",
X"03E8",
X"055F",
X"0271",
X"FB9B",
X"FAA1",
X"FE89",
X"04E2",
X"04E2",
X"03E8",
X"FC18",
X"FAA1",
X"FD12",
X"0465",
X"055F",
X"01F4",
X"FAA1",
X"FB1E",
X"FC18",
X"036B",
X"055F",
X"036B",
X"FC18",
X"FAA1",
X"FD12",
X"0465",
X"055F",
X"01F4",
X"FB1E",
X"FB9B",
X"FB9B",
X"036B",
X"055F",
X"036B",
X"FC18",
X"FAA1",
X"FD8F",
X"04E2",
X"04E2",
X"0271",
X"FB1E",
X"FAA1",
X"FB9B",
X"0465",
X"05DC",
X"02EE",
X"FB9B",
X"FA24",
X"FD8F",
X"04E2",
X"04E2",
X"0465",
X"FC95",
X"FAA1",
X"FC95",
X"03E8",
X"05DC",
X"0271",
X"FB9B",
X"FA24",
X"FE0C",
X"055F",
X"055F",
X"0465",
X"FB9B",
X"FA24",
X"FD12",
X"0465",
X"05DC",
X"0271",
X"FAA1",
X"FAA1",
X"FB9B",
X"036B",
X"05DC",
X"036B",
X"FC18",
X"F9A7",
X"FD12",
X"0465",
X"05DC",
X"01F4",
X"FAA1",
X"FAA1",
X"FB9B",
X"03E8",
X"05DC",
X"036B",
X"FB9B",
X"FA24",
X"FD12",
X"055F",
X"055F",
X"0465",
X"FC95",
X"F9A7",
X"FC95",
X"03E8",
X"05DC",
X"02EE",
X"FB9B",
X"F9A7",
X"FD8F",
X"055F",
X"055F",
X"0465",
X"FC95",
X"FA24",
X"FC95",
X"03E8",
X"05DC",
X"036B",
X"FB1E",
X"FA24",
X"FB9B",
X"036B",
X"05DC",
X"03E8",
X"FC18",
X"FA24",
X"FC95",
X"0465",
X"0659",
X"02EE",
X"FAA1",
X"FAA1",
X"FB9B",
X"02EE",
X"05DC",
X"03E8",
X"FC95",
X"FA24",
X"FC95",
X"0465",
X"05DC",
X"036B",
X"FB1E",
X"FA24",
X"FB1E",
X"036B",
X"0659",
X"03E8",
X"FC18",
X"F9A7",
X"FC95",
X"04E2",
X"055F",
X"04E2",
X"FD12",
X"FA24",
X"FC18",
X"02EE",
X"0659",
X"03E8",
X"FC18",
X"F9A7",
X"FC95",
X"04E2",
X"055F",
X"055F",
X"FC95",
X"F9A7",
X"FB9B",
X"03E8",
X"0659",
X"03E8",
X"FB9B",
X"FAA1",
X"FAA1",
X"0271",
X"05DC",
X"0465",
X"FD12",
X"F9A7",
X"FB9B",
X"036B",
X"05DC",
X"036B",
X"FB9B",
X"FAA1",
X"FAA1",
X"0271",
X"05DC",
X"0465",
X"FD12",
X"FA24",
X"FB9B",
X"0465",
X"055F",
X"055F",
X"FE0C",
X"F9A7",
X"FB1E",
X"0271",
X"05DC",
X"0465",
X"FD12",
X"F9A7",
X"FC18",
X"0465",
X"055F",
X"055F",
X"FE0C",
X"FA24",
X"FB1E",
X"0271",
X"05DC",
X"0465",
X"FC95",
X"FA24",
X"FB1E",
X"0271",
X"055F",
X"04E2",
X"FE0C",
X"FA24",
X"FB9B",
X"02EE",
X"05DC",
X"03E8",
X"FC18",
X"FB1E",
X"FAA1",
X"0177",
X"05DC",
X"04E2",
X"FE0C",
X"FA24",
X"FB9B",
X"0271",
X"055F",
X"0465",
X"FC18",
X"FAA1",
X"FAA1",
X"0177",
X"05DC",
X"04E2",
X"FD8F",
X"FA24",
X"FB9B",
X"036B",
X"04E2",
X"055F",
X"FE89",
X"FAA1",
X"FB1E",
X"0177",
X"055F",
X"04E2",
X"FD12",
X"FAA1",
X"FC18",
X"036B",
X"04E2",
X"055F",
X"FE89",
X"FAA1",
X"FB1E",
X"0271",
X"05DC",
X"0465",
X"FC95",
X"FB1E",
X"FAA1",
X"007D",
X"04E2",
X"04E2",
X"FE89",
X"FA24",
X"FB9B",
X"0271",
X"05DC",
X"03E8",
X"FC95",
X"FB1E",
X"FAA1",
X"00FA",
X"055F",
X"04E2",
X"FE0C",
X"FAA1",
X"FB1E",
X"02EE",
X"055F",
X"04E2",
X"FF83",
X"FAA1",
X"FB1E",
X"0177",
X"05DC",
X"0465",
X"FE0C",
X"FA24",
X"FB9B",
X"02EE",
X"04E2",
X"055F",
X"FF83",
X"FAA1",
X"FB1E",
X"0177",
X"055F",
X"04E2",
X"FE0C",
X"FB1E",
X"FB9B",
X"0271",
X"055F",
X"055F",
X"FF06",
X"FAA1",
X"FB1E",
X"01F4",
X"055F",
X"0465",
X"FD12",
X"FAA1",
X"FAA1",
X"0000",
X"055F",
X"04E2",
X"FE89",
X"FAA1",
X"FB1E",
X"01F4",
X"05DC",
X"04E2",
X"FD12",
X"FB1E",
X"FAA1",
X"007D",
X"05DC",
X"055F",
X"FE89",
X"FA24",
X"FAA1",
X"0271",
X"055F",
X"05DC",
X"FF83",
X"FAA1",
X"FAA1",
X"00FA",
X"05DC",
X"055F",
X"FE0C",
X"FA24",
X"FB1E",
X"0271",
X"055F",
X"055F",
X"FF83",
X"FA24",
X"FAA1",
X"0177",
X"0659",
X"05DC",
X"FD8F",
X"FA24",
X"FAA1",
X"0000",
X"05DC",
X"055F",
X"FF06",
X"F9A7",
X"FB1E",
X"0177",
X"0659",
X"04E2",
X"FD12",
X"FAA1",
X"FA24",
X"0000",
X"05DC",
X"055F",
X"FF06",
X"F9A7",
X"FAA1",
X"01F4",
X"05DC",
X"055F",
X"0000",
X"FAA1",
X"FB1E",
X"007D",
X"05DC",
X"04E2",
X"FE89",
X"FA24",
X"FB1E",
X"01F4",
X"055F",
X"055F",
X"007D",
X"FAA1",
X"FB1E",
X"007D",
X"055F",
X"04E2",
X"FE89",
X"FAA1",
X"FB1E",
X"01F4",
X"055F",
X"055F",
X"0000",
X"FAA1",
X"FB1E",
X"00FA",
X"055F",
X"04E2",
X"FE89",
X"FAA1",
X"FAA1",
X"FF06",
X"055F",
X"055F",
X"FF83",
X"FAA1",
X"FB1E",
X"00FA",
X"055F",
X"04E2",
X"FE0C",
X"FB1E",
X"FAA1",
X"FF83",
X"055F",
X"055F",
X"FF83",
X"FAA1",
X"FAA1",
X"00FA",
X"055F",
X"055F",
X"00FA",
X"FB1E",
X"FAA1",
X"FF83",
X"055F",
X"04E2",
X"FF83",
X"FAA1",
X"FB1E",
X"0177",
X"04E2",
X"04E2",
X"00FA",
X"FAA1",
X"FAA1",
X"0000",
X"055F",
X"055F",
X"FF06",
X"FAA1",
X"FB1E",
X"FE89",
X"055F",
X"055F",
X"007D",
X"FAA1",
X"FB1E",
X"0000",
X"055F",
X"04E2",
X"FF06",
X"FB1E",
X"FAA1",
X"FE89",
X"055F",
X"055F",
X"007D",
X"FA24",
X"FAA1",
X"007D",
X"055F",
X"05DC",
X"0177",
X"FAA1",
X"FAA1",
X"FF06",
X"055F",
X"055F",
X"0000",
X"FAA1",
X"FAA1",
X"007D",
X"055F",
X"055F",
X"01F4",
X"FAA1",
X"FAA1",
X"FF06",
X"055F",
X"055F",
X"007D",
X"FB1E",
X"FA24",
X"007D",
X"055F",
X"055F",
X"0177",
X"FAA1",
X"FA24",
X"FF83",
X"055F",
X"05DC",
X"0000",
X"FAA1",
X"FAA1",
X"FE0C",
X"04E2",
X"055F",
X"0177",
X"FB1E",
X"FAA1",
X"FF83",
X"055F",
X"05DC",
X"FF83",
X"FAA1",
X"FAA1",
X"FE0C",
X"04E2",
X"05DC",
X"00FA",
X"FB1E",
X"FAA1",
X"FF83",
X"055F",
X"055F",
X"0271",
X"FB1E",
X"FAA1",
X"FE0C",
X"055F",
X"055F",
X"00FA",
X"FB1E",
X"FAA1",
X"0000",
X"055F",
X"055F",
X"0271",
X"FB1E",
X"FAA1",
X"FE89",
X"04E2",
X"05DC",
X"007D",
X"FAA1",
X"FB1E",
X"FD12",
X"04E2",
X"055F",
X"01F4",
X"FB1E",
X"FAA1",
X"FE89",
X"04E2",
X"055F",
X"007D",
X"FB1E",
X"FB1E",
X"FD12",
X"0465",
X"055F",
X"01F4",
X"FB1E",
X"FAA1",
X"FF06",
X"04E2",
X"055F",
X"0271",
X"FB9B",
X"FB1E",
X"FE0C",
X"0465",
X"055F",
X"0177",
X"FB9B",
X"FB1E",
X"FF06",
X"04E2",
X"04E2",
X"02EE",
X"FB9B",
X"FB1E",
X"FE0C",
X"03E8",
X"04E2",
X"0177",
X"FB9B",
X"FAA1",
X"FF83",
X"04E2",
X"04E2",
X"0271",
X"FB9B",
X"FAA1",
X"FE0C",
X"0465",
X"055F",
X"00FA",
X"FB1E",
X"FB1E",
X"FD12",
X"0465",
X"04E2",
X"0271",
X"FB9B",
X"FAA1",
X"FE89",
X"0465",
X"055F",
X"007D",
X"FB1E",
X"FB1E",
X"FD12",
X"0465",
X"055F",
X"0271",
X"FB9B",
X"FAA1",
X"FE89",
X"04E2",
X"04E2",
X"036B",
X"FC18",
X"FAA1",
X"FD12",
X"0465",
X"055F",
X"01F4",
X"FB9B",
X"FAA1",
X"FF06",
X"04E2",
X"04E2",
X"02EE",
X"FC18",
X"FAA1",
X"FD8F",
X"0465",
X"05DC",
X"01F4",
X"FAA1",
X"FB1E",
X"FC95",
X"03E8",
X"055F",
X"02EE",
X"FC18",
X"FAA1",
X"FE0C",
X"0465",
X"055F",
X"0177",
X"FB1E",
X"FB1E",
X"FC95",
X"03E8",
X"055F",
X"0271",
X"FB9B",
X"FAA1",
X"FE0C",
X"04E2",
X"04E2",
X"01F4",
X"FB1E",
X"FAA1",
X"FC95",
X"03E8",
X"05DC",
X"01F4",
X"FB9B",
X"FAA1",
X"FE0C",
X"055F",
X"04E2",
X"036B",
X"FC18",
X"FAA1",
X"FD12",
X"03E8",
X"055F",
X"01F4",
X"FB9B",
X"FAA1",
X"FE89",
X"04E2",
X"04E2",
X"036B",
X"FC18",
X"FA24",
X"FD8F",
X"0465",
X"055F",
X"01F4",
X"FB1E",
X"FB1E",
X"FC95",
X"036B",
X"04E2",
X"036B",
X"FC95",
X"FAA1",
X"FE0C",
X"03E8",
X"055F",
X"0177",
X"FB1E",
X"FB1E",
X"FC18",
X"036B",
X"055F",
X"02EE",
X"FB9B",
X"FAA1",
X"FD8F",
X"04E2",
X"0465",
X"03E8",
X"FD12",
X"FAA1",
X"FC95",
X"036B",
X"055F",
X"0271",
X"FC18",
X"FAA1",
X"FE0C",
X"04E2",
X"04E2",
X"03E8",
X"FD12",
X"FAA1",
X"FC95",
X"03E8",
X"055F",
X"0271",
X"FB1E",
X"FB1E",
X"FC18",
X"036B",
X"055F",
X"036B",
X"FC95",
X"FAA1",
X"FD8F",
X"03E8",
X"055F",
X"0271",
X"FB9B",
X"FB9B",
X"FC18",
X"02EE",
X"055F",
X"036B",
X"FC95",
X"FB1E",
X"FD8F",
X"03E8",
X"04E2",
X"0271",
X"FB9B",
X"FB1E",
X"FC18",
X"02EE",
X"055F",
X"02EE",
X"FC95",
X"FB1E",
X"FD8F",
X"0465",
X"0465",
X"03E8",
X"FD12",
X"FB1E",
X"FC95",
X"02EE",
X"055F",
X"02EE",
X"FC95",
X"FAA1",
X"FD8F",
X"0465",
X"0465",
X"0465",
X"FD12",
X"FB1E",
X"FC95",
X"036B",
X"04E2",
X"0271",
X"FC18",
X"FB9B",
X"FC18",
X"0271",
X"04E2",
X"036B",
X"FD8F",
X"FB1E",
X"FD12",
X"02EE",
X"04E2",
X"0271",
X"FC18",
X"FB9B",
X"FC18",
X"0271",
X"04E2",
X"036B",
X"FD12",
X"FB1E",
X"FD12",
X"03E8",
X"03E8",
X"03E8",
X"FE0C",
X"FB1E",
X"FC95",
X"0271",
X"04E2",
X"02EE",
X"FD12",
X"FB9B",
X"FD12",
X"03E8",
X"0465",
X"03E8",
X"FE0C",
X"FB1E",
X"FC95",
X"02EE",
X"04E2",
X"02EE",
X"FC95",
X"FB9B",
X"FC18",
X"01F4",
X"0465",
X"036B",
X"FD8F",
X"FB1E",
X"FD12",
X"02EE",
X"0465",
X"02EE",
X"FC95",
X"FB9B",
X"FB9B",
X"01F4",
X"04E2",
X"036B",
X"FD8F",
X"FB1E",
X"FD12",
X"02EE",
X"04E2",
X"02EE",
X"FC95",
X"FB1E",
X"FB9B",
X"01F4",
X"055F",
X"036B",
X"FD12",
X"FB1E",
X"FC95",
X"036B",
X"0465",
X"0465",
X"FE0C",
X"FAA1",
X"FC18",
X"01F4",
X"04E2",
X"036B",
X"FD8F",
X"FB1E",
X"FC95",
X"036B",
X"0465",
X"0465",
X"FE0C",
X"FAA1",
X"FC18",
X"0271",
X"04E2",
X"036B",
X"FD12",
X"FB9B",
X"FB9B",
X"0177",
X"055F",
X"03E8",
X"FE0C",
X"FAA1",
X"FC18",
X"0271",
X"04E2",
X"036B",
X"FC95",
X"FB9B",
X"FB1E",
X"0177",
X"04E2",
X"0465",
X"FD8F",
X"FB1E",
X"FC18",
X"02EE",
X"0465",
X"0465",
X"FF06",
X"FAA1",
X"FC18",
X"01F4",
X"055F",
X"03E8",
X"FD8F",
X"FB9B",
X"FC95",
X"02EE",
X"0465",
X"04E2",
X"FE89",
X"FB1E",
X"FC18",
X"01F4",
X"04E2",
X"03E8",
X"FD8F",
X"FB9B",
X"FB9B",
X"0177",
X"0465",
X"03E8",
X"FE89",
X"FB1E",
X"FC95",
X"01F4",
X"0465",
X"036B",
X"FD12",
X"FC18",
X"FB9B",
X"00FA",
X"04E2",
X"03E8",
X"FE89",
X"FB9B",
X"FC95",
X"01F4",
X"0465",
X"036B",
X"FD12",
X"FB9B",
X"FB9B",
X"00FA",
X"04E2",
X"03E8",
X"FE0C",
X"FB9B",
X"FC95",
X"0271",
X"0465",
X"0465",
X"FF83",
X"FB1E",
X"FC18",
X"00FA",
X"0465",
X"036B",
X"FE0C",
X"FB1E",
X"FC95",
X"02EE",
X"03E8",
X"0465",
X"FF06",
X"FB1E",
X"FC18",
X"01F4",
X"04E2",
X"036B",
X"FD8F",
X"FB9B",
X"FB9B",
X"007D",
X"04E2",
X"0465",
X"FF06",
X"FB1E",
X"FC18",
X"01F4",
X"04E2",
X"03E8",
X"FD8F",
X"FB9B",
X"FB1E",
X"007D",
X"0465",
X"0465",
X"FF06",
X"FB1E",
X"FB9B",
X"01F4",
X"0465",
X"0465",
X"0000",
X"FB9B",
X"FB9B",
X"007D",
X"04E2",
X"0465",
X"FF06",
X"FB9B",
X"FC18",
X"01F4",
X"0465",
X"04E2",
X"0000",
X"FB9B",
X"FB9B",
X"0000",
X"0465",
X"0465",
X"FF06",
X"FB9B",
X"FB1E",
X"0000",
X"0465",
X"04E2",
X"0000",
X"FB9B",
X"FB9B",
X"007D",
X"0465",
X"0465",
X"FE89",
X"FB9B",
X"FB1E",
X"FF83",
X"0465",
X"0465",
X"0000",
X"FB9B",
X"FB9B",
X"007D",
X"04E2",
X"0465",
X"FE89",
X"FB1E",
X"FB1E",
X"FF83",
X"04E2",
X"04E2",
X"FF83",
X"FB1E",
X"FB9B",
X"0177",
X"04E2",
X"0465",
X"007D",
X"FB1E",
X"FB9B",
X"FF83",
X"0465",
X"0465",
X"FF06",
X"FB1E",
X"FB9B",
X"01F4",
X"0465",
X"04E2",
X"007D",
X"FB1E",
X"FB1E",
X"007D",
X"0465",
X"0465",
X"FE89",
X"FB9B",
X"FB9B",
X"FF06",
X"0465",
X"04E2",
X"007D",
X"FB1E",
X"FB9B",
X"00FA",
X"04E2",
X"0465",
X"FE89",
X"FB9B",
X"FB9B",
X"FF83",
X"0465",
X"0465",
X"0000",
X"FB9B",
X"FB9B",
X"00FA",
X"0465",
X"0465",
X"00FA",
X"FB9B",
X"FB9B",
X"FF83",
X"0465",
X"03E8",
X"FF83",
X"FB9B",
X"FC18",
X"0177",
X"0465",
X"0465",
X"00FA",
X"FB9B",
X"FC18",
X"FF83",
X"0465",
X"0465",
X"FF83",
X"FB9B",
X"FB9B",
X"007D",
X"0465",
X"0465",
X"007D",
X"FB9B",
X"FB9B",
X"0000",
X"0465",
X"0465",
X"FF06",
X"FB9B",
X"FB9B",
X"FE89",
X"0465",
X"0465",
X"007D",
X"FB9B",
X"FB9B",
X"0000",
X"04E2",
X"0465",
X"FF06",
X"FB9B",
X"FB9B",
X"FF06",
X"0465",
X"0465",
X"0000",
X"FB9B",
X"FB9B",
X"007D",
X"0465",
X"0465",
X"0177",
X"FB9B",
X"FB9B",
X"FF06",
X"0465",
X"04E2",
X"0000",
X"FB1E",
X"FB9B",
X"00FA",
X"0465",
X"0465",
X"0177",
X"FB9B",
X"FB9B",
X"FF83",
X"0465",
X"0465",
X"0000",
X"FB9B",
X"FB9B",
X"FE0C",
X"0465",
X"04E2",
X"0177",
X"FB9B",
X"FB9B",
X"0000",
X"04E2",
X"0465",
X"FF83",
X"FB9B",
X"FB9B",
X"FE89",
X"0465",
X"0465",
X"00FA",
X"FB9B",
X"FB1E",
X"FF83",
X"0465",
X"04E2",
X"01F4",
X"FC18",
X"FB9B",
X"FE89",
X"0465",
X"0465",
X"007D",
X"FB9B",
X"FB1E",
X"0000",
X"0465",
X"0465",
X"01F4",
X"FC18",
X"FB9B",
X"FE89",
X"03E8",
X"04E2",
X"007D",
X"FC18",
X"FB1E",
X"FF83",
X"0465",
X"04E2",
X"01F4",
X"FB9B",
X"FB1E",
X"FE89",
X"03E8",
X"04E2",
X"007D",
X"FB9B",
X"FB9B",
X"FD8F",
X"03E8",
X"0465",
X"0177",
X"FC95",
X"FB1E",
X"FF06",
X"0465",
X"04E2",
X"0000",
X"FB9B",
X"FC18",
X"FE0C",
X"03E8",
X"0465",
X"0177",
X"FC18",
X"FB1E",
X"FF06",
X"0465",
X"0465",
X"02EE",
X"FC95",
X"FB9B",
X"FE0C",
X"03E8",
X"04E2",
X"0177",
X"FB9B",
X"FB1E",
X"FF83",
X"0465",
X"03E8",
X"0271",
X"FC95",
X"FB9B",
X"FE0C",
X"036B",
X"0465",
X"00FA",
X"FB9B",
X"FB9B",
X"FC95",
X"036B",
X"0465",
X"01F4",
X"FC95",
X"FB1E",
X"FE89",
X"03E8",
X"04E2",
X"00FA",
X"FC18",
X"FC18",
X"FD8F",
X"036B",
X"0465",
X"01F4",
X"FC95",
X"FB9B",
X"FE89",
X"03E8",
X"0465",
X"02EE",
X"FC95",
X"FB9B",
X"FD8F",
X"02EE",
X"0465",
X"01F4",
X"FC95",
X"FB9B",
X"FF06",
X"03E8",
X"03E8",
X"02EE",
X"FC95",
X"FB9B",
X"FE0C",
X"02EE",
X"0465",
X"0177",
X"FC95",
X"FB9B",
X"FF06",
X"03E8",
X"03E8",
X"02EE",
X"FC95",
X"FB9B",
X"FE0C",
X"036B",
X"0465",
X"0177",
X"FC95",
X"FC18",
X"FD12",
X"02EE",
X"0465",
X"01F4",
X"FD12",
X"FB9B",
X"FE89",
X"03E8",
X"0465",
X"00FA",
X"FC18",
X"FC95",
X"FD8F",
X"02EE",
X"0465",
X"01F4",
X"FC95",
X"FB9B",
X"FE89",
X"03E8",
X"03E8",
X"036B",
X"FD12",
X"FB9B",
X"FD8F",
X"036B",
X"04E2",
X"0177",
X"FC18",
X"FB9B",
X"FF06",
X"03E8",
X"03E8",
X"02EE",
X"FD12",
X"FB9B",
X"FE0C",
X"036B",
X"0465",
X"0177",
X"FC18",
X"FC95",
X"FD12",
X"02EE",
X"0465",
X"01F4",
X"FC95",
X"FB9B",
X"FE89",
X"036B",
X"0465",
X"00FA",
X"FB9B",
X"FC95",
X"FD8F",
X"036B",
X"03E8",
X"01F4",
X"FC95",
X"FC18",
X"FE89",
X"03E8",
X"03E8",
X"0271",
X"FD12",
X"FC18",
X"FD8F",
X"02EE",
X"03E8",
X"0177",
X"FD12",
X"FC18",
X"FE89",
X"03E8",
X"03E8",
X"02EE",
X"FD12",
X"FB9B",
X"FE0C",
X"02EE",
X"03E8",
X"0177",
X"FC95",
X"FC18",
X"FE89",
X"03E8",
X"036B",
X"02EE",
X"FD8F",
X"FC18",
X"FD8F",
X"02EE",
X"03E8",
X"01F4",
X"FC95",
X"FC18",
X"FC95",
X"0271",
X"0465",
X"02EE",
X"FD8F",
X"FB9B",
X"FE0C",
X"036B",
X"0465",
X"01F4",
X"FC18",
X"FC18",
X"FC95",
X"01F4",
X"03E8",
X"02EE",
X"FD12",
X"FC18",
X"FD8F",
X"036B",
X"03E8",
X"03E8",
X"FE0C",
X"FB9B",
X"FC95",
X"0271",
X"0465",
X"0271",
X"FD12",
X"FB9B",
X"FE0C",
X"036B",
X"03E8",
X"036B",
X"FD8F",
X"FB9B",
X"FD12",
X"0271",
X"0465",
X"0271",
X"FC95",
X"FC95",
X"FC18",
X"0177",
X"0465",
X"02EE",
X"FE0C",
X"FB9B",
X"FD8F",
X"0271",
X"0465",
X"0271",
X"FC95",
X"FC18",
X"FC95",
X"01F4",
X"0465",
X"02EE",
X"FD8F",
X"FB9B",
X"FD8F",
X"02EE",
X"03E8",
X"0271",
X"FD12",
X"FC18",
X"FC95",
X"01F4",
X"0465",
X"02EE",
X"FD8F",
X"FB9B",
X"FD12",
X"02EE",
X"03E8",
X"03E8",
X"FE0C",
X"FB9B",
X"FD12",
X"01F4",
X"0465",
X"02EE",
X"FD8F",
X"FB9B",
X"FD8F",
X"036B",
X"036B",
X"036B",
X"FE0C",
X"FC18",
X"FD12",
X"0271",
X"0465",
X"0271",
X"FD12",
X"FC18",
X"FC95",
X"01F4",
X"0465",
X"036B",
X"FE0C",
X"FB9B",
X"FD12",
X"02EE",
X"0465",
X"0271",
X"FC95",
X"FC18",
X"FC95",
X"01F4",
X"0465",
X"02EE",
X"FD8F",
X"FB9B",
X"FD12",
X"036B",
X"03E8",
X"036B",
X"FE89",
X"FB9B",
X"FC95",
X"01F4",
X"0465",
X"02EE",
X"FD8F",
X"FB9B",
X"FD12",
X"036B",
X"03E8",
X"036B",
X"FE0C",
X"FB9B",
X"FD12",
X"0271",
X"0465",
X"02EE",
X"FD12",
X"FC18",
X"FC95",
X"0177",
X"0465",
X"036B",
X"FE0C",
X"FB9B",
X"FD12",
X"01F4",
X"03E8",
X"02EE",
X"FD12",
X"FC18",
X"FC18",
X"0177",
X"0465",
X"02EE",
X"FE0C",
X"FC18",
X"FD12",
X"0271",
X"0465",
X"02EE",
X"FD12",
X"FC18",
X"FC18",
X"0177",
X"0465",
X"036B",
X"FE0C",
X"FB9B",
X"FC95",
X"0271",
X"03E8",
X"03E8",
X"FF06",
X"FB9B",
X"FC95",
X"0177",
X"0465",
X"036B",
X"FE0C",
X"FC18",
X"FD12",
X"02EE",
X"03E8",
X"03E8",
X"FF06",
X"FC18",
X"FC95",
X"01F4",
X"0465",
X"036B",
X"FD8F",
X"FC18",
X"FC95",
X"007D",
X"0465",
X"03E8",
X"FE89",
X"FB9B",
X"FC95",
X"01F4",
X"0465",
X"02EE",
X"FD8F",
X"FC18",
X"FC18",
X"00FA",
X"0465",
X"03E8",
X"FE89",
X"FB9B",
X"FC95",
X"0271",
X"03E8",
X"03E8",
X"FF83",
X"FB9B",
X"FC18",
X"00FA",
X"0465",
X"036B",
X"FE89",
X"FB9B",
X"FC95",
X"0271",
X"03E8",
X"0465",
X"FF83",
X"FB9B",
X"FC18",
X"00FA",
X"0465",
X"03E8",
X"FE0C",
X"FB9B",
X"FC18",
X"007D",
X"03E8",
X"03E8",
X"FF06",
X"FC18",
X"FC18",
X"0177",
X"03E8",
X"03E8",
X"FE0C",
X"FC18",
X"FC18",
X"0000",
X"0465",
X"03E8",
X"FF06",
X"FC18",
X"FC18",
X"00FA",
X"0465",
X"036B",
X"FE0C",
X"FC18",
X"FB9B",
X"007D",
X"0465",
X"03E8",
X"FF06",
X"FB9B",
X"FC18",
X"0177",
X"03E8",
X"03E8",
X"007D",
X"FC18",
X"FC18",
X"007D",
X"03E8",
X"03E8",
X"FF06",
X"FC18",
X"FC95",
X"01F4",
X"03E8",
X"03E8",
X"0000",
X"FC18",
X"FC18",
X"007D",
X"03E8",
X"03E8",
X"FE89",
X"FC18",
X"FC95",
X"FF83",
X"036B",
X"036B",
X"FF83",
X"FC95",
X"FC18",
X"007D",
X"03E8",
X"036B",
X"FE89",
X"FC95",
X"FC18",
X"FF83",
X"036B",
X"036B",
X"FF83",
X"FC18",
X"FC95",
X"0177",
X"036B",
X"03E8",
X"007D",
X"FC18",
X"FC95",
X"007D",
X"03E8",
X"036B",
X"FF83",
X"FC18",
X"FC95",
X"0177",
X"036B",
X"036B",
X"007D",
X"FC18",
X"FC95",
X"007D",
X"03E8",
X"036B",
X"FF06",
X"FC18",
X"FC95",
X"0000",
X"036B",
X"036B",
X"FF83",
X"FC95",
X"FD12",
X"00FA",
X"036B",
X"036B",
X"FE89",
X"FC18",
X"FD12",
X"FF83",
X"03E8",
X"02EE",
X"FF83",
X"FC18",
X"FC95",
X"007D",
X"03E8",
X"02EE",
X"FE89",
X"FC95",
X"FC95",
X"0000",
X"03E8",
X"036B",
X"FF83",
X"FC18",
X"FC95",
X"00FA",
X"03E8",
X"02EE",
X"007D",
X"FC95",
X"FD12",
X"0000",
X"036B",
X"036B",
X"FF06",
X"FC95",
X"FD12",
X"0177",
X"03E8",
X"02EE",
X"007D",
X"FC95",
X"FC95",
X"007D",
X"03E8",
X"02EE",
X"FF06",
X"FC18",
X"FD12",
X"FF06",
X"036B",
X"036B",
X"0000",
X"FC95",
X"FC95",
X"007D",
X"036B",
X"02EE",
X"FF06",
X"FC95",
X"FC95",
X"FF83",
X"036B",
X"036B",
X"0000",
X"FC95",
X"FC95",
X"007D",
X"036B",
X"036B",
X"00FA",
X"FC95",
X"FC95",
X"FF83",
X"036B",
X"036B",
X"0000",
X"FC95",
X"FC18",
X"007D",
X"036B",
X"036B",
X"00FA",
X"FC95",
X"FC95",
X"FF83",
X"036B",
X"03E8",
X"0000",
X"FC18",
X"FC95",
X"FF06",
X"036B",
X"036B",
X"00FA",
X"FC95",
X"FC95",
X"FF83",
X"036B",
X"036B",
X"0000",
X"FC18",
X"FC95",
X"FE89",
X"036B",
X"036B",
X"00FA",
X"FC95",
X"FC18",
X"FF83",
X"036B",
X"03E8",
X"0000",
X"FC18",
X"FC95",
X"FE89",
X"03E8",
X"03E8",
X"007D",
X"FC18",
X"FC18",
X"0000",
X"03E8",
X"03E8",
X"01F4",
X"FC95",
X"FC18",
X"FF06",
X"036B",
X"03E8",
X"007D",
X"FC95",
X"FC18",
X"0000",
X"03E8",
X"03E8",
X"0177",
X"FC95",
X"FB9B",
X"FF06",
X"03E8",
X"03E8",
X"007D",
X"FC18",
X"FC18",
X"FE0C",
X"036B",
X"0465",
X"0177",
X"FC95",
X"FB9B",
X"FF06",
X"036B",
X"0465",
X"007D",
X"FC18",
X"FC18",
X"FE0C",
X"036B",
X"0465",
X"0177",
X"FC95",
X"FB9B",
X"FF06",
X"03E8",
X"03E8",
X"0271",
X"FC95",
X"FC18",
X"FE89",
X"036B",
X"0465",
X"00FA",
X"FD12",
X"FB9B",
X"FF83",
X"03E8",
X"03E8",
X"01F4",
X"FC95",
X"FC18",
X"FE89",
X"02EE",
X"03E8",
X"00FA",
X"FC95",
X"FC18",
X"FF06",
X"036B",
X"03E8",
X"01F4",
X"FC95",
X"FC18",
X"FE89",
X"036B",
X"03E8",
X"00FA",
X"FC95",
X"FC95",
X"FE0C",
X"02EE",
X"03E8",
X"0177",
X"FD12",
X"FC18",
X"FE89",
X"036B",
X"03E8",
X"007D",
X"FC18",
X"FC95",
X"FD8F",
X"036B",
X"03E8",
X"0177",
X"FC95",
X"FC18",
X"FF06",
X"036B",
X"036B",
X"0271",
X"FD12",
X"FC18",
X"FE0C",
X"02EE",
X"03E8",
X"0177",
X"FD12",
X"FC18",
X"FF06",
X"036B",
X"036B",
X"0271",
X"FD12",
X"FC18",
X"FE89",
X"02EE",
X"03E8",
X"0177",
X"FC95",
X"FC95",
X"FD12",
X"0271",
X"03E8",
X"01F4",
X"FD12",
X"FC18",
X"FE89",
X"02EE",
X"03E8",
X"00FA",
X"FC95",
X"FC95",
X"FD8F",
X"02EE",
X"03E8",
X"01F4",
X"FD8F",
X"FC18",
X"FE89",
X"036B",
X"036B",
X"02EE",
X"FD8F",
X"FC18",
X"FD8F",
X"0271",
X"03E8",
X"01F4",
X"FD8F",
X"FC18",
X"FE89",
X"02EE",
X"02EE",
X"02EE",
X"FD8F",
X"FC95",
X"FE0C",
X"0271",
X"036B",
X"01F4",
X"FD12",
X"FC95",
X"FE89",
X"036B",
X"036B",
X"02EE",
X"FD8F",
X"FC18",
X"FD8F",
X"02EE",
X"03E8",
X"0177",
X"FD12",
X"FC95",
X"FD12",
X"0271",
X"03E8",
X"0271",
X"FD8F",
X"FC18",
X"FE0C",
X"0271",
X"03E8",
X"0177",
X"FC95",
X"FC95",
X"FD12",
X"0271",
X"03E8",
X"01F4",
X"FD12",
X"FC18",
X"FE89",
X"02EE",
X"036B",
X"02EE",
X"FE0C",
X"FC18",
X"FD8F",
X"0271",
X"03E8",
X"01F4",
X"FD8F",
X"FC95",
X"FE89",
X"02EE",
X"036B",
X"02EE",
X"FE0C",
X"FC18",
X"FD8F",
X"0271",
X"036B",
X"01F4",
X"FD12",
X"FD12",
X"FD12",
X"01F4",
X"03E8",
X"0271",
X"FE0C",
X"FC18",
X"FE0C",
X"0271",
X"036B",
X"01F4",
X"FD12",
X"FD12",
X"FD12",
X"01F4",
X"036B",
X"0271",
X"FE0C",
X"FC95",
X"FE0C",
X"0271",
X"036B",
X"02EE",
X"FE0C",
X"FD12",
X"FD8F",
X"01F4",
X"036B",
X"01F4",
X"FE0C",
X"FC95",
X"FE0C",
X"02EE",
X"02EE",
X"02EE",
X"FE89",
X"FC95",
X"FD8F",
X"01F4",
X"036B",
X"01F4",
X"FE0C",
X"FC95",
X"FE0C",
X"02EE",
X"02EE",
X"02EE",
X"FE0C",
X"FC95",
X"FD8F",
X"01F4",
X"036B",
X"01F4",
X"FD8F",
X"FD12",
X"FD12",
X"0177",
X"036B",
X"0271",
X"FE89",
X"FC95",
X"FD8F",
X"01F4",
X"036B",
X"01F4",
X"FD8F",
X"FD12",
X"FD12",
X"0177",
X"036B",
X"0271",
X"FE0C",
X"FC95",
X"FD8F",
X"0271",
X"02EE",
X"02EE",
X"FE89",
X"FC95",
X"FD8F",
X"0177",
X"03E8",
X"0271",
X"FE0C",
X"FC95",
X"FD8F",
X"0271",
X"036B",
X"036B",
X"FE89",
X"FC95",
X"FD12",
X"01F4",
X"03E8",
X"0271",
X"FD8F",
X"FC95",
X"FC95",
X"00FA",
X"03E8",
X"02EE",
X"FE89",
X"FC95",
X"FD8F",
X"01F4",
X"036B",
X"0271",
X"FD8F",
X"FC95",
X"FC95",
X"0177",
X"036B",
X"02EE",
X"FE89",
X"FC95",
X"FD12",
X"01F4",
X"036B",
X"036B",
X"FE89",
X"FC95",
X"FD12",
X"0177",
X"036B",
X"0271",
X"FE89",
X"FC95",
X"FD8F",
X"0271",
X"02EE",
X"036B",
X"FF06",
X"FC95",
X"FD12",
X"0177",
X"036B",
X"0271",
X"FE89",
X"FC95",
X"FD12",
X"0271",
X"036B",
X"036B",
X"FF06",
X"FC95",
X"FD12",
X"0177",
X"036B",
X"02EE",
X"FE0C",
X"FD12",
X"FC95",
X"007D",
X"036B",
X"02EE",
X"FF06",
X"FC95",
X"FD8F",
X"0177",
X"036B",
X"0271",
X"FE0C",
X"FD12",
X"FC95",
X"00FA",
X"036B",
X"02EE",
X"FE89",
X"FC95",
X"FD8F",
X"0177",
X"02EE",
X"036B",
X"FF83",
X"FC95",
X"FD12",
X"00FA",
X"036B",
X"0271",
X"FE89",
X"FD12",
X"FD8F",
X"0177",
X"02EE",
X"036B",
X"FF83",
X"FD12",
X"FD12",
X"00FA",
X"02EE",
X"02EE",
X"FE89",
X"FD12",
X"FC95",
X"007D",
X"02EE",
X"02EE",
X"FF06",
X"FD12",
X"FD8F",
X"00FA",
X"02EE",
X"0271",
X"FE89",
X"FD12",
X"FD12",
X"007D",
X"02EE",
X"02EE",
X"FF06",
X"FD12",
X"FD8F",
X"00FA",
X"02EE",
X"02EE",
X"FE89",
X"FD12",
X"FD12",
X"007D",
X"036B",
X"0271",
X"FF06",
X"FC95",
X"FD8F",
X"0177",
X"02EE",
X"02EE",
X"FF83",
X"FD12",
X"FD12",
X"007D",
X"036B",
X"0271",
X"FF06",
X"FD12",
X"FD12",
X"01F4",
X"02EE",
X"02EE",
X"FF83",
X"FC95",
X"FD12",
X"00FA",
X"036B",
X"02EE",
X"FE89",
X"FD12",
X"FC95",
X"0000",
X"036B",
X"02EE",
X"FF83",
X"FC95",
X"FD12",
X"00FA",
X"036B",
X"02EE",
X"FE89",
X"FD12",
X"FC95",
X"0000",
X"036B",
X"036B",
X"FF83",
X"FC95",
X"FD12",
X"0177",
X"036B",
X"036B",
X"0000",
X"FC95",
X"FD12",
X"007D",
X"036B",
X"02EE",
X"FF06",
X"FC95",
X"FD12",
X"0177",
X"02EE",
X"036B",
X"0000",
X"FC95",
X"FC95",
X"007D",
X"036B",
X"02EE",
X"FE89",
X"FC95",
X"FC95",
X"0000",
X"036B",
X"02EE",
X"FF83",
X"FD12",
X"FD12",
X"00FA",
X"036B",
X"02EE",
X"FE89",
X"FD12",
X"FD12",
X"0000",
X"02EE",
X"02EE",
X"FF83",
X"FD12",
X"FD12",
X"00FA",
X"02EE",
X"02EE",
X"FF06",
X"FD12",
X"FD12",
X"0000",
X"036B",
X"02EE",
X"FF83",
X"FC95",
X"FD12",
X"0177",
X"02EE",
X"02EE",
X"007D",
X"FD12",
X"FD12",
X"0000",
X"02EE",
X"02EE",
X"FF83",
X"FD12",
X"FD12",
X"00FA",
X"02EE",
X"02EE",
X"007D",
X"FD12",
X"FD12",
X"0000",
X"02EE",
X"02EE",
X"FF06",
X"FD12",
X"FD12",
X"FF83",
X"02EE",
X"02EE",
X"0000",
X"FD12",
X"FD12",
X"007D",
X"02EE",
X"02EE",
X"FF06",
X"FD12",
X"FC95",
X"FF83",
X"02EE",
X"02EE",
X"0000",
X"FD12",
X"FD12",
X"007D",
X"02EE",
X"02EE",
X"00FA",
X"FD12",
X"FD12",
X"FF83",
X"02EE",
X"02EE",
X"FF83",
X"FD12",
X"FD12",
X"007D",
X"02EE",
X"02EE",
X"007D",
X"FD12",
X"FD12",
X"0000",
X"02EE",
X"02EE",
X"FF83",
X"FD12",
X"FD12",
X"FF06",
X"0271",
X"02EE",
X"007D",
X"FD8F",
X"FD12",
X"0000",
X"02EE",
X"02EE",
X"FF83",
X"FD12",
X"FD8F",
X"FF06",
X"0271",
X"02EE",
X"007D",
X"FD8F",
X"FD8F",
X"0000",
X"0271",
X"0271",
X"0000",
X"FD12",
X"FD12",
X"FF06",
X"02EE",
X"0271",
X"0000",
X"FD8F",
X"FD12",
X"007D",
X"02EE",
X"0271",
X"00FA",
X"FD8F",
X"FD12",
X"FF83",
X"0271",
X"02EE",
X"0000",
X"FD8F",
X"FD12",
X"007D",
X"02EE",
X"0271",
X"00FA",
X"FD8F",
X"FD12",
X"FF83",
X"0271",
X"02EE",
X"0000",
X"FD12",
X"FD8F",
X"FE89",
X"0271",
X"02EE",
X"00FA",
X"FD8F",
X"FD12",
X"0000",
X"02EE",
X"02EE",
X"FF83",
X"FD12",
X"FD12",
X"FF06",
X"0271",
X"02EE",
X"007D",
X"FD12",
X"FD12",
X"0000",
X"02EE",
X"02EE",
X"0177",
X"FD8F",
X"FD12",
X"FF06",
X"0271",
X"02EE",
X"007D",
X"FD8F",
X"FD12",
X"0000",
X"02EE",
X"02EE",
X"0177",
X"FD8F",
X"FD12",
X"FF83",
X"02EE",
X"02EE",
X"007D",
X"FD12",
X"FD12",
X"FE89",
X"0271",
X"02EE",
X"00FA",
X"FD8F",
X"FD12",
X"FF83",
X"0271",
X"02EE",
X"007D",
X"FD12",
X"FD12",
X"FE89",
X"0271",
X"036B",
X"00FA",
X"FD8F",
X"FD12",
X"FF06",
X"0271",
X"02EE",
X"007D",
X"FD12",
X"FD12",
X"FE89",
X"0271",
X"02EE",
X"00FA",
X"FD8F",
X"FD12",
X"FF83",
X"02EE",
X"02EE",
X"01F4",
X"FD8F",
X"FC95",
X"FE89",
X"0271",
X"036B",
X"00FA",
X"FD12",
X"FD12",
X"FF83",
X"02EE",
X"02EE",
X"0177",
X"FD8F",
X"FD12",
X"FF06",
X"0271",
X"02EE",
X"007D",
X"FD12",
X"FD12",
X"FE0C",
X"0271",
X"02EE",
X"0177",
X"FD8F",
X"FC95",
X"FF06",
X"02EE",
X"02EE",
X"007D",
X"FD12",
X"FD12",
X"FE89",
X"0271",
X"02EE",
X"00FA",
X"FD8F",
X"FD12",
X"FF83",
X"02EE",
X"0271",
X"01F4",
X"FE0C",
X"FD12",
X"FE89",
X"0271",
X"02EE",
X"00FA",
X"FD8F",
X"FD12",
X"FF83",
X"02EE",
X"0271",
X"01F4",
X"FD8F",
X"FD12",
X"FE89",
X"0271",
X"02EE",
X"00FA",
X"FD8F",
X"FD8F",
X"FE89",
X"0271",
X"0271",
X"0177",
X"FD8F",
X"FD12",
X"FF06",
X"0271",
X"02EE",
X"00FA",
X"FD12",
X"FD8F",
X"FE0C",
X"01F4",
X"02EE",
X"0177",
X"FD8F",
X"FD12",
X"FF06",
X"0271",
X"02EE",
X"00FA",
X"FD8F",
X"FD8F",
X"FE89",
X"01F4",
X"02EE",
X"0177",
X"FE0C",
X"FD12",
X"FF06",
X"0271",
X"0271",
X"01F4",
X"FE0C",
X"FD12",
X"FE89",
X"01F4",
X"02EE",
X"0177",
X"FD8F",
X"FD12",
X"FF06",
X"0271",
X"0271",
X"01F4",
X"FE0C",
X"FD12",
X"FE89",
X"01F4",
X"02EE",
X"0177",
X"FD8F",
X"FD8F",
X"FD8F",
X"0177",
X"02EE",
X"01F4",
X"FE0C",
X"FD12",
X"FE89",
X"01F4",
X"02EE",
X"00FA",
X"FD8F",
X"FD8F",
X"FE0C",
X"0177",
X"02EE",
X"01F4",
X"FE0C",
X"FD12",
X"FE89",
X"0271",
X"0271",
X"0271",
X"FE89",
X"FD12",
X"FE0C",
X"01F4",
X"02EE",
X"0177",
X"FE0C",
X"FD12",
X"FE89",
X"0271",
X"0271",
X"0271",
X"FE89",
X"FD12",
X"FE0C",
X"01F4",
X"02EE",
X"0177",
X"FE0C",
X"FD8F",
X"FE89",
X"0271",
X"02EE",
X"01F4",
X"FE0C",
X"FD8F",
X"FE89",
X"01F4",
X"0271",
X"0177",
X"FD8F",
X"FD8F",
X"FD8F",
X"0177",
X"02EE",
X"0177",
X"FE0C",
X"FD12",
X"FE89",
X"01F4",
X"02EE",
X"00FA",
X"FD8F",
X"FD8F",
X"FE0C",
X"01F4",
X"0271",
X"0177",
X"FE0C",
X"FD8F",
X"FE89",
X"0271",
X"0271",
X"01F4",
X"FE89",
X"FD8F",
X"FE89",
X"0177",
X"02EE",
X"0177",
X"FE0C",
X"FD12",
X"FF06",
X"0271",
X"0271",
X"01F4",
X"FE89",
X"FD8F",
X"FE89",
X"01F4",
X"0271",
X"0177",
X"FD8F",
X"FE0C",
X"FE0C",
X"00FA",
X"0271",
X"01F4",
X"FE89",
X"FD8F",
X"FE89",
X"01F4",
X"0271",
X"0177",
X"FD8F",
X"FD8F",
X"FE0C",
X"0177",
X"0271",
X"0177",
X"FE0C",
X"FD8F",
X"FE89",
X"01F4",
X"0271",
X"01F4",
X"FF06",
X"FD8F",
X"FE89",
X"0177",
X"0271",
X"0177",
X"FE89",
X"FD8F",
X"FE89",
X"0271",
X"0271",
X"01F4",
X"FF06",
X"FD8F",
X"FE89",
X"0177",
X"0271",
X"0177",
X"FE0C",
X"FD8F",
X"FE89",
X"01F4",
X"0271",
X"01F4",
X"FE89",
X"FD8F",
X"FE0C",
X"0177",
X"0271",
X"0177",
X"FE0C",
X"FD8F",
X"FE0C",
X"00FA",
X"0271",
X"01F4",
X"FE89",
X"FD12",
X"FE0C",
X"0177",
X"02EE",
X"0177",
X"FD8F",
X"FD8F",
X"FE0C",
X"0177",
X"0271",
X"01F4",
X"FE89",
X"FD8F",
X"FE89",
X"01F4",
X"0271",
X"0271",
X"FF06",
X"FD8F",
X"FE0C",
X"00FA",
X"02EE",
X"01F4",
X"FE89",
X"FD12",
X"FE0C",
X"01F4",
X"0271",
X"01F4",
X"FF06",
X"FD8F",
X"FE0C",
X"0177",
X"0271",
X"01F4",
X"FE89",
X"FD8F",
X"FD8F",
X"007D",
X"0271",
X"01F4",
X"FF06",
X"FD8F",
X"FE0C",
X"00FA",
X"0271",
X"01F4",
X"FE89",
X"FD8F",
X"FD8F",
X"007D",
X"0271",
X"01F4",
X"FF06",
X"FD8F",
X"FE0C",
X"0177",
X"0271",
X"0271",
X"FF83",
X"FD8F",
X"FE0C",
X"007D",
X"0271",
X"01F4",
X"FF06",
X"FD8F",
X"FE0C",
X"0177",
X"0271",
X"0271",
X"FF83",
X"FD8F",
X"FE0C",
X"00FA",
X"0271",
X"01F4",
X"FF06",
X"FD8F",
X"FE0C",
X"0177",
X"01F4",
X"0271",
X"FF83",
X"FD8F",
X"FE0C",
X"00FA",
X"0271",
X"01F4",
X"FF06",
X"FE0C",
X"FD8F",
X"0000",
X"0271",
X"01F4",
X"FF83",
X"FD8F",
X"FE0C",
X"00FA",
X"0271",
X"01F4",
X"FE89",
X"FE0C",
X"FD8F",
X"007D",
X"0271",
X"01F4",
X"FF83",
X"FD8F",
X"FE0C",
X"00FA",
X"01F4",
X"0271",
X"0000",
X"FD8F",
X"FD8F",
X"007D",
X"0271",
X"01F4",
X"FF83",
X"FD8F",
X"FE0C",
X"00FA",
X"01F4",
X"0271",
X"0000",
X"FD8F",
X"FE0C",
X"007D",
X"0271",
X"01F4",
X"FF06",
X"FE0C",
X"FD8F",
X"FF83",
X"0271",
X"0271",
X"0000",
X"FD8F",
X"FD8F",
X"007D",
X"0271",
X"01F4",
X"FF06",
X"FE0C",
X"FD8F",
X"0000",
X"0271",
X"0271",
X"FF83",
X"FD8F",
X"FD8F",
X"00FA",
X"0271",
X"01F4",
X"0000",
X"FE0C",
X"FD8F",
X"0000",
X"0271",
X"01F4",
X"FF83",
X"FD8F",
X"FE0C",
X"00FA",
X"01F4",
X"0271",
X"007D",
X"FD8F",
X"FD8F",
X"0000",
X"0271",
X"01F4",
X"FF83",
X"FD8F",
X"FE0C",
X"00FA",
X"01F4",
X"0271",
X"0000",
X"FD8F",
X"FE0C",
X"007D",
X"0271",
X"01F4",
X"FF06",
X"FD8F",
X"FD8F",
X"0000",
X"0271",
X"0271",
X"0000",
X"FD8F",
X"FE0C",
X"007D",
X"0271",
X"01F4",
X"FF06",
X"FD8F",
X"FD8F",
X"0000",
X"0271",
X"01F4",
X"FF83",
X"FD8F",
X"FE0C",
X"007D",
X"0271",
X"0271",
X"007D",
X"FD8F",
X"FD8F",
X"0000",
X"0271",
X"01F4",
X"FF83",
X"FD8F",
X"FE0C",
X"00FA",
X"01F4",
X"01F4",
X"0000",
X"FE0C",
X"FE0C",
X"0000",
X"0271",
X"01F4",
X"FF83",
X"FE0C",
X"FE0C",
X"FF83",
X"01F4",
X"01F4",
X"0000",
X"FE0C",
X"FD8F",
X"007D",
X"0271",
X"01F4",
X"FF06",
X"FE0C",
X"FE0C",
X"FF83",
X"01F4",
X"0271",
X"0000",
X"FD8F",
X"FE0C",
X"007D",
X"0271",
X"01F4",
X"FF83",
X"FE0C",
X"FD8F",
X"FF83",
X"0271",
X"0271",
X"0000",
X"FE0C",
X"FD8F",
X"007D",
X"01F4",
X"0271",
X"00FA",
X"FE0C",
X"FD8F",
X"FF83",
X"0271",
X"0271",
X"0000",
X"FE0C",
X"FD8F",
X"007D",
X"01F4",
X"01F4",
X"007D",
X"FE0C",
X"FD8F",
X"0000",
X"01F4",
X"0271",
X"0000",
X"FE0C",
X"FD8F",
X"FF06",
X"01F4",
X"0271",
X"007D",
X"FE0C",
X"FD8F",
X"0000",
X"01F4",
X"0271",
X"FF83",
X"FE0C",
X"FD8F",
X"FF83",
X"01F4",
X"0271",
X"0000",
X"FE0C",
X"FE0C",
X"0000",
X"0271",
X"01F4",
X"00FA",
X"FE0C",
X"FD8F",
X"FF83",
X"0271",
X"0271",
X"0000",
X"FD8F",
X"FD8F",
X"007D",
X"0271",
X"01F4",
X"00FA",
X"FE0C",
X"FD8F",
X"FF83",
X"0271",
X"0271",
X"0000",
X"FE0C",
X"FE0C",
X"FF06",
X"01F4",
X"0271",
X"007D",
X"FE0C",
X"FD8F",
X"FF83",
X"0271",
X"0271",
X"0000",
X"FD8F",
X"FE0C",
X"FF06",
X"01F4",
X"0271",
X"007D",
X"FE0C",
X"FD8F",
X"0000",
X"0271",
X"01F4",
X"0000",
X"FE0C",
X"FD8F",
X"FF06",
X"01F4",
X"0271",
X"007D",
X"FE0C",
X"FD8F",
X"0000",
X"0271",
X"01F4",
X"00FA",
X"FE0C",
X"FD8F",
X"FF83",
X"01F4",
X"0271",
X"0000",
X"FE0C",
X"FD8F",
X"0000",
X"0271",
X"01F4",
X"00FA",
X"FE0C",
X"FD8F",
X"FF83",
X"01F4",
X"0271",
X"007D",
X"FD8F",
X"FE0C",
X"FF06",
X"01F4",
X"0271",
X"007D",
X"FE0C",
X"FD8F",
X"FF83",
X"01F4",
X"0271",
X"0000",
X"FE0C",
X"FE0C",
X"FF06",
X"01F4",
X"0271",
X"007D",
X"FE0C",
X"FE0C",
X"FF83",
X"01F4",
X"01F4",
X"0177",
X"FE0C",
X"FD8F",
X"FF06",
X"01F4",
X"01F4",
X"007D",
X"FE0C",
X"FE0C",
X"0000",
X"01F4",
X"01F4",
X"00FA",
X"FE89",
X"FE0C",
X"FF06",
X"01F4",
X"0271",
X"007D",
X"FE0C",
X"FE0C",
X"FE89",
X"0177",
X"01F4",
X"00FA",
X"FE89",
X"FE0C",
X"FF06",
X"01F4",
X"01F4",
X"007D",
X"FE0C",
X"FE0C",
X"FE89",
X"0177",
X"01F4",
X"00FA",
X"FE89",
X"FE0C",
X"FF83",
X"01F4",
X"01F4",
X"007D",
X"FE0C",
X"FE0C",
X"FF06",
X"0177",
X"01F4",
X"00FA",
X"FE89",
X"FE0C",
X"FF83",
X"01F4",
X"01F4",
X"0177",
X"FE89",
X"FE0C",
X"FF06",
X"0177",
X"01F4",
X"007D",
X"FE0C",
X"FE0C",
X"FF83",
X"01F4",
X"01F4",
X"0177",
X"FE89",
X"FE0C",
X"FF06",
X"0177",
X"0271",
X"00FA",
X"FE0C",
X"FE0C",
X"FE89",
X"0177",
X"01F4",
X"00FA",
X"FE89",
X"FE0C",
X"FF06",
X"0177",
X"01F4",
X"007D",
X"FE0C",
X"FE0C",
X"FE89",
X"0177",
X"01F4",
X"00FA",
X"FE89",
X"FE0C",
X"FF06",
X"01F4",
X"01F4",
X"0177",
X"FE89",
X"FE0C",
X"FE89",
X"0177",
X"01F4",
X"00FA",
X"FE89",
X"FE0C",
X"FF83",
X"01F4",
X"01F4",
X"0177",
X"FE89",
X"FE0C",
X"FF06",
X"0177",
X"0271",
X"00FA",
X"FE0C",
X"FE0C",
X"FE89",
X"0177",
X"01F4",
X"0177",
X"FE89",
X"FE0C",
X"FF06",
X"0177",
X"01F4",
X"00FA",
X"FE0C",
X"FE0C",
X"FE89",
X"0177",
X"01F4",
X"0177",
X"FE89",
X"FE0C",
X"FF06",
X"0177",
X"01F4",
X"00FA",
X"FE89",
X"FE0C",
X"FE89",
X"00FA",
X"01F4",
X"0177",
X"FE89",
X"FE0C",
X"FF06",
X"0177",
X"01F4",
X"01F4",
X"FF06",
X"FE0C",
X"FE89",
X"0177",
X"01F4",
X"00FA",
X"FE89",
X"FE0C",
X"FF06",
X"01F4",
X"01F4",
X"0177",
X"FF06",
X"FE0C",
X"FE89",
X"0177",
X"01F4",
X"0177",
X"FE89",
X"FE0C",
X"FE0C",
X"00FA",
X"01F4",
X"0177",
X"FE89",
X"FE0C",
X"FF06",
X"0177",
X"01F4",
X"00FA",
X"FE89",
X"FE0C",
X"FE89",
X"00FA",
X"01F4",
X"0177",
X"FE89",
X"FE0C",
X"FF06",
X"0177",
X"01F4",
X"01F4",
X"FF06",
X"FE0C",
X"FE89",
X"00FA",
X"01F4",
X"00FA",
X"FE89",
X"FE0C",
X"FF06",
X"0177",
X"01F4",
X"0177",
X"FF06",
X"FE0C",
X"FE89",
X"0177",
X"01F4",
X"00FA",
X"FE89",
X"FE0C",
X"FE89",
X"00FA",
X"0177",
X"0177",
X"FF06",
X"FE0C",
X"FF06",
X"00FA",
X"01F4",
X"00FA",
X"FE89",
X"FE89",
X"FE89",
X"00FA",
X"01F4",
X"0177",
X"FF06",
X"FE0C",
X"FF06",
X"00FA",
X"01F4",
X"00FA",
X"FE89",
X"FE89",
X"FE89",
X"00FA",
X"01F4",
X"0177",
X"FF06",
X"FE0C",
X"FF06",
X"0177",
X"0177",
X"0177",
X"FF06",
X"FE0C",
X"FE89",
X"00FA",
X"01F4",
X"00FA",
X"FF06",
X"FE0C",
X"FF06",
X"0177",
X"0177",
X"0177",
X"FF06",
X"FE0C",
X"FE89",
X"00FA",
X"01F4",
X"00FA",
X"FE89",
X"FE89",
X"FE89",
X"007D",
X"01F4",
X"0177",
X"FF06",
X"FE0C",
X"FF06",
X"0177",
X"01F4",
X"00FA",
X"FE89",
X"FE89",
X"FE89",
X"00FA",
X"01F4",
X"0177",
X"FF06",
X"FE0C",
X"FF06",
X"0177",
X"0177",
X"0177",
X"FF83",
X"FE0C",
X"FE89",
X"00FA",
X"01F4",
X"0177",
X"FF06",
X"FE0C",
X"FF06",
X"0177",
X"01F4",
X"0177",
X"FF83",
X"FE0C",
X"FE89",
X"00FA",
X"01F4",
X"0177",
X"FF06",
X"FE0C",
X"FE89",
X"0177",
X"01F4",
X"0177",
X"FF06",
X"FE0C",
X"FE89",
X"00FA",
X"01F4",
X"0177",
X"FE89",
X"FE0C",
X"FE0C",
X"007D",
X"01F4",
X"0177",
X"FF06",
X"FE0C",
X"FE89",
X"00FA",
X"01F4",
X"0177",
X"FE89",
X"FE0C",
X"FE89",
X"007D",
X"01F4",
X"0177",
X"FF06",
X"FE0C",
X"FE89",
X"00FA",
X"01F4",
X"01F4",
X"FF83",
X"FE0C",
X"FE0C",
X"007D",
X"01F4",
X"0177",
X"FF06",
X"FE0C",
X"FE89",
X"0177",
X"01F4",
X"0177",
X"FF83",
X"FE0C",
X"FE89",
X"00FA",
X"01F4",
X"0177",
X"FF06",
X"FE0C",
X"FE89",
X"0000",
X"01F4",
X"01F4",
X"FF83",
X"FE0C",
X"FE89",
X"00FA",
X"01F4",
X"0177",
X"FF06",
X"FE89",
X"FE0C",
X"007D",
X"01F4",
X"01F4",
X"FF83",
X"FE0C",
X"FE89",
X"00FA",
X"01F4",
X"01F4",
X"0000",
X"FE0C",
X"FE89",
X"007D",
X"01F4",
X"0177",
X"FF83",
X"FE0C",
X"FE89",
X"00FA",
X"0177",
X"0177",
X"0000",
X"FE0C",
X"FE89",
X"007D",
X"0177",
X"0177",
X"FF83",
X"FE89",
X"FE89",
X"00FA",
X"01F4",
X"01F4",
X"0000",
X"FE0C",
X"FE89",
X"007D",
X"01F4",
X"0177",
X"FF83",
X"FE89",
X"FE89",
X"0000",
X"01F4",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"007D",
X"0177",
X"0177",
X"FF06",
X"FE89",
X"FE89",
X"0000",
X"01F4",
X"0177",
X"FF83",
X"FE89",
X"FE89",
X"007D",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE0C",
X"0000",
X"01F4",
X"0177",
X"FF83",
X"FE89",
X"FE89",
X"007D",
X"0177",
X"01F4",
X"0000",
X"FE89",
X"FE0C",
X"0000",
X"0177",
X"0177",
X"FF83",
X"FE89",
X"FE89",
X"FF83",
X"0177",
X"01F4",
X"0000",
X"FE89",
X"FE89",
X"007D",
X"0177",
X"0177",
X"FF83",
X"FE89",
X"FE0C",
X"0000",
X"01F4",
X"01F4",
X"0000",
X"FE89",
X"FE0C",
X"007D",
X"01F4",
X"01F4",
X"0000",
X"FE89",
X"FE0C",
X"0000",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"007D",
X"0177",
X"0177",
X"007D",
X"FE89",
X"FE89",
X"0000",
X"0177",
X"0177",
X"FF83",
X"FE89",
X"FE89",
X"007D",
X"0177",
X"0177",
X"0000",
X"FE0C",
X"FE89",
X"0000",
X"0177",
X"0177",
X"FF83",
X"FE89",
X"FE89",
X"FF83",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"0000",
X"0177",
X"0177",
X"FF83",
X"FE89",
X"FE89",
X"FF83",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"0000",
X"0177",
X"0177",
X"007D",
X"FE89",
X"FE89",
X"0000",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"007D",
X"0177",
X"0177",
X"007D",
X"FE89",
X"FE89",
X"0000",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"FF83",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"0000",
X"0177",
X"0177",
X"FF83",
X"FE89",
X"FE89",
X"FF83",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"0000",
X"0177",
X"0177",
X"007D",
X"FE89",
X"FE89",
X"FF83",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"0000",
X"0177",
X"0177",
X"007D",
X"FE89",
X"FE89",
X"0000",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"0000",
X"0177",
X"0177",
X"007D",
X"FE89",
X"FE89",
X"0000",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"FF83",
X"0177",
X"0177",
X"007D",
X"FF06",
X"FE89",
X"0000",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"FF83",
X"0177",
X"0177",
X"007D",
X"FE89",
X"FE89",
X"0000",
X"0177",
X"0177",
X"007D",
X"FE89",
X"FE89",
X"FF83",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"0000",
X"0177",
X"0177",
X"007D",
X"FE89",
X"FE89",
X"FF83",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"FF06",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FE89",
X"FF83",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"FF06",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FE89",
X"FF83",
X"00FA",
X"0177",
X"007D",
X"FE89",
X"FE89",
X"FF83",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FE89",
X"FF83",
X"0177",
X"00FA",
X"00FA",
X"FF06",
X"FE89",
X"FF83",
X"00FA",
X"0177",
X"007D",
X"FE89",
X"FE89",
X"0000",
X"0177",
X"00FA",
X"007D",
X"FF06",
X"FE89",
X"FF83",
X"0177",
X"0177",
X"0000",
X"FE89",
X"FE89",
X"FF06",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FE89",
X"FF83",
X"0177",
X"00FA",
X"0000",
X"FE89",
X"FF06",
X"FF83",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FF06",
X"0000",
X"0177",
X"00FA",
X"00FA",
X"FF06",
X"FE89",
X"FF83",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FE89",
X"0000",
X"0177",
X"00FA",
X"007D",
X"FF06",
X"FE89",
X"FF83",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FF06",
X"FF06",
X"00FA",
X"00FA",
X"007D",
X"FF06",
X"FF06",
X"FF83",
X"00FA",
X"00FA",
X"007D",
X"FF06",
X"FF06",
X"FF06",
X"00FA",
X"00FA",
X"007D",
X"FF06",
X"FF06",
X"FF83",
X"00FA",
X"00FA",
X"007D",
X"FF06",
X"FF06",
X"FF06",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FE89",
X"FF83",
X"00FA",
X"00FA",
X"00FA",
X"FF06",
X"FE89",
X"FF83",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FE89",
X"FF83",
X"00FA",
X"00FA",
X"00FA",
X"FF06",
X"FE89",
X"FF06",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FF06",
X"FF06",
X"00FA",
X"0177",
X"00FA",
X"FF06",
X"FE89",
X"FF83",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FF06",
X"FF06",
X"00FA",
X"0177",
X"00FA",
X"FF06",
X"FE89",
X"FF83",
X"00FA",
X"00FA",
X"00FA",
X"FF06",
X"FE89",
X"FF06",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FE89",
X"FF83",
X"00FA",
X"00FA",
X"00FA",
X"FF06",
X"FE89",
X"FF06",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF06",
X"FE89",
X"FF83",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FF06",
X"FF06",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FE89",
X"FF83",
X"00FA",
X"00FA",
X"007D",
X"FF06",
X"FF06",
X"FF06",
X"007D",
X"0177",
X"00FA",
X"FF06",
X"FE89",
X"FF83",
X"00FA",
X"00FA",
X"00FA",
X"FF83",
X"FE89",
X"FF06",
X"007D",
X"00FA",
X"007D",
X"FF06",
X"FF06",
X"FF83",
X"00FA",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"007D",
X"FF06",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"007D",
X"FF06",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"00FA",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF83",
X"00FA",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"00FA",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"007D",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"FF83",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"00FA",
X"00FA",
X"0000",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF06",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"0000",
X"0000",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"0000",
X"0000",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"FF83",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D"





 );

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
      if (ENA='1') then
		Q_tmp <= sin_table(conv_integer(ADDR));
--		if conv_integer(ADDR) < 6294 then
--		   Done <= '1';
--		end if;	
		else 
		 Q_tmp <= ( others => '0');
      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end arch;